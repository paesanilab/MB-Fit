netcdf x2b_A1B2Z2_D1E2_v1x {
  // global attributes 
  :name = "x2b_A1B2Z2_D1E2_v1x<3>";
  :d_intra_AB =  9.456180336306371e-01; // A^(-1))
  :k_intra_AB =  1.012210945112919e+00; // A^(-1))
  :d_intra_BB =  1.478734942157645e-01; // A^(-1))
  :k_intra_BB =  8.687447666922434e-01; // A^(-1))
  :d_intra_DE =  1.562363345817676e+00; // A^(-1))
  :k_intra_DE =  1.178074665863358e+00; // A^(-1))
  :d_intra_EE =  5.833090049789817e-01; // A^(-1))
  :k_intra_EE =  1.817125247843581e+00; // A^(-1))
  :d_AD =  9.368104072408366e-02; // A^(-1))
  :k_AD =  1.967402295403801e+00; // A^(-1))
  :d_AE =  8.054394432416823e-01; // A^(-1))
  :k_AE =  2.974430053069379e+00; // A^(-1))
  :d_BD =  6.271199705824921e+00; // A^(-1))
  :k_BD =  9.014396154830446e-01; // A^(-1))
  :d_BE =  6.726600251761202e+00; // A^(-1))
  :k_BE =  1.673367133446074e+00; // A^(-1))
  :d_DZ =  2.087864453786822e+00; // A^(-1))
  :k_DZ =  1.435959164515135e+00; // A^(-1))
  :d_EZ =  4.045839071180502e+00; // A^(-1))
  :k_EZ =  2.058738367691483e+00; // A^(-1))
  :r2i =  6.000000000000000e+00; // A
  :r2f =  7.000000000000000e+00; // A
  dimensions:
  poly = 492;
  variables:
    double poly(poly);
data:
poly =
 4.692249405592280e-02, // 0
-1.739055794173007e+02, // 1
-5.905311757265770e+02, // 2
-1.343068207498834e+00, // 3
 8.496413525246860e-01, // 4
-2.979098286875208e+01, // 5
-1.344830018629170e-02, // 6
-6.202570916604831e+00, // 7
 2.314406363814029e+00, // 8
-5.703881588175485e+02, // 9
 4.323153921986059e+00, // 10
-3.478985551806785e+01, // 11
-1.412095768313563e+03, // 12
 1.657917006316609e+02, // 13
-4.264168427137235e-02, // 14
 1.589119532185932e+00, // 15
-4.260718741836011e-01, // 16
-6.995347623217705e-04, // 17
 7.441953977407140e+00, // 18
 2.607654106315471e-05, // 19
 2.024924432714684e+00, // 20
 5.467379158365636e+01, // 21
-1.068889252281304e-05, // 22
-5.876992805950923e-04, // 23
-3.881828216881688e-06, // 24
-8.729325156275873e+02, // 25
 3.061310060607843e+03, // 26
-5.892288066144836e-01, // 27
 2.324935055043330e-02, // 28
-3.229075065723959e+02, // 29
 2.146312937088803e+02, // 30
 9.378201251612757e-07, // 31
-1.729286086745818e+00, // 32
-4.738652200604655e-05, // 33
 1.438781220488233e-02, // 34
-1.880002925457927e-02, // 35
 6.581268653733072e-03, // 36
-4.441130506718799e-02, // 37
 6.715681173054625e+00, // 38
-4.191384542784913e-02, // 39
 1.399279418395447e-01, // 40
-3.454810064698524e-07, // 41
 2.439144870997241e+00, // 42
-4.018696795293526e+01, // 43
-4.801678914806155e+02, // 44
-8.817068961677319e+01, // 45
 2.012940169988176e+03, // 46
-1.376027920328277e+03, // 47
-1.863512791744055e-01, // 48
 1.253682418980304e+03, // 49
 9.481226227637611e+02, // 50
 2.686172988438295e-01, // 51
-3.764520967531124e+02, // 52
 3.697963164359584e-02, // 53
-8.293473863080605e+02, // 54
-1.644484342902469e-02, // 55
 6.062221484518963e-07, // 56
 6.960724722562066e-01, // 57
 2.580684921440745e+03, // 58
-3.597193844694480e-02, // 59
 1.097078474576679e+02, // 60
 1.489637921703165e+00, // 61
-3.152070434641033e+00, // 62
 3.079913118482489e+00, // 63
 3.251218378175150e-02, // 64
 1.228082702738589e+03, // 65
-1.181572663133814e+03, // 66
-5.642014070320004e+02, // 67
 3.601366663011046e+03, // 68
 7.155718050864389e-02, // 69
-3.375492102116772e-08, // 70
 1.648473857446126e-04, // 71
-3.353358594987348e-03, // 72
-7.796637781496895e-01, // 73
 5.603756996719955e-02, // 74
 1.211600561607447e-04, // 75
-1.329268654090868e-06, // 76
-2.322671022950957e+03, // 77
-7.183739680022403e+01, // 78
-1.818227186024918e-03, // 79
-2.596147937639139e+00, // 80
-6.128193321118743e-07, // 81
 6.046277365207786e-06, // 82
 1.138710273069088e-04, // 83
 6.612013846811000e-03, // 84
 1.057174097856002e+01, // 85
 3.456014202424046e-03, // 86
-1.774441012167662e+02, // 87
-1.425308916369667e+01, // 88
-7.212758680270496e+02, // 89
-2.856477779242534e+01, // 90
 6.685094319186173e+01, // 91
-1.484449557135822e+03, // 92
 8.923749033266925e-07, // 93
 1.681401686746638e-04, // 94
-1.865437324941834e+01, // 95
-4.473832092984711e-02, // 96
 3.861215597565261e-01, // 97
-1.462959558793381e-03, // 98
 1.384875475922984e-01, // 99
-1.087063189645135e+02, // 100
 5.828043472014290e-02, // 101
 6.578137294199532e+02, // 102
-1.316679792692027e+01, // 103
-3.733028652037943e-11, // 104
-2.202908135388299e-01, // 105
 4.830400273392295e-03, // 106
 1.313615559529967e-06, // 107
 4.148382367383633e-05, // 108
 2.798041785134196e+00, // 109
 8.374914022796038e-08, // 110
 1.052334373747879e-01, // 111
 2.611116909688923e-03, // 112
 5.408115765315169e-06, // 113
-2.554278445854690e-05, // 114
 4.636070819254758e-01, // 115
 4.378186944138699e-06, // 116
 7.902187098314342e-01, // 117
 1.439794406171961e+01, // 118
-9.807253777234196e-04, // 119
 1.663780148841081e+01, // 120
-1.845908524576441e-08, // 121
 7.138928713617191e-05, // 122
 3.754573883587038e-04, // 123
-4.115474618600982e-05, // 124
-1.436671696651808e+02, // 125
 9.347040755739179e-02, // 126
-7.162926485463317e-02, // 127
 2.772261211704630e-02, // 128
-8.811505913036742e-01, // 129
 2.414922987333426e+03, // 130
-3.800486991006388e-04, // 131
-7.676785834122313e-01, // 132
-4.357150369097537e+03, // 133
-9.396916393716053e+02, // 134
-1.378209430861691e+02, // 135
-6.383744641671008e+00, // 136
 3.396580902439786e-03, // 137
-2.502842795691950e-01, // 138
-4.010864128021546e-05, // 139
-9.310741227622126e+00, // 140
-2.419379804471994e-04, // 141
-2.410238413027779e+01, // 142
 1.148421566668836e-05, // 143
-4.992303861981693e-05, // 144
 1.847503147404503e-10, // 145
 2.251308989689271e-01, // 146
-1.576094657573316e-01, // 147
-1.226008484227842e-02, // 148
 1.393668206424080e-04, // 149
-5.137301406855380e-03, // 150
 6.470621942791197e-04, // 151
 1.511721173063983e-05, // 152
-2.493659532115139e-03, // 153
-1.067666750972777e-07, // 154
-8.020378446564046e-04, // 155
 1.153128644787601e+02, // 156
-1.260536461336939e+00, // 157
 2.624374206115509e+01, // 158
-3.151286809782675e-04, // 159
 1.048705865456938e+01, // 160
-1.054966963479851e+03, // 161
-4.855095598126230e-04, // 162
-1.568091961555292e+01, // 163
 9.036056255541800e-03, // 164
-1.573022855355932e-04, // 165
-4.739573582624839e-05, // 166
 1.892180366071654e-06, // 167
 8.126840054321796e+00, // 168
-1.778064228927384e+03, // 169
 3.694907344518451e-03, // 170
-5.011367584775326e-07, // 171
-2.611648785954328e-02, // 172
-3.790132903478045e-06, // 173
-6.287728550428940e-06, // 174
 3.747938401828057e-06, // 175
 3.507235158968478e-02, // 176
 6.667832234065882e-03, // 177
 4.047265725222470e-09, // 178
-4.420485533266151e+00, // 179
 3.755944005329472e-05, // 180
-5.962434072113932e+02, // 181
-9.537379662988877e-01, // 182
 9.404488660887203e+02, // 183
-1.956232332979731e+00, // 184
-5.010320512734613e+02, // 185
 4.013922261268398e-02, // 186
 1.389122189001417e-07, // 187
-3.123241233787739e-09, // 188
-2.788043846625130e+00, // 189
 3.833669595925114e-04, // 190
-3.288743388612309e+00, // 191
 2.665184643885212e+01, // 192
-1.411729322391187e+00, // 193
 6.146329452228021e-03, // 194
-4.190292880141714e-03, // 195
-3.341876606599329e-07, // 196
 1.822612505001294e-07, // 197
 1.560214342412246e-06, // 198
 1.182434840423064e-03, // 199
-7.081697827366741e+02, // 200
-7.700699607916544e-09, // 201
-1.227897089136872e-04, // 202
 2.847610241681447e-05, // 203
 6.261965605237045e-02, // 204
-1.094375014000638e-02, // 205
-8.677414398812072e-03, // 206
 4.457129360617781e-01, // 207
-1.023900655104266e+00, // 208
-7.272390792329031e-01, // 209
-9.532935390994346e-08, // 210
-7.566413084898066e+00, // 211
-9.557797980024096e+02, // 212
 2.565351608343845e+00, // 213
-5.566710681173690e-05, // 214
 1.345213166035974e-02, // 215
-2.109408976322957e-03, // 216
-5.068376639399649e-02, // 217
-5.049828597124481e-03, // 218
 1.001259321648540e+02, // 219
 6.882200177787261e+01, // 220
 2.101121894355265e-01, // 221
 8.245667954817607e-07, // 222
 4.533532932644166e-03, // 223
-1.960977156358575e+00, // 224
-4.051442641951956e-07, // 225
-2.689469988113346e-08, // 226
-4.729243241489798e+02, // 227
 4.265745757402863e-05, // 228
 2.888262249066528e-01, // 229
-1.969705628804270e+03, // 230
 1.595279955347539e-01, // 231
 1.615451396854343e-04, // 232
 8.836637348573759e-02, // 233
-6.935801798034434e-02, // 234
 4.354949677731248e+01, // 235
-2.343092474588791e-02, // 236
-9.965042612026540e-02, // 237
-2.876335191334131e+02, // 238
 1.722302377410664e+01, // 239
 9.826514920282756e-03, // 240
 9.770370102841151e-07, // 241
-2.092260285892473e+02, // 242
-6.357765213938789e-05, // 243
 7.527556106599357e-07, // 244
-2.721072132210338e-09, // 245
-2.972480737142288e-01, // 246
-4.860913552460889e+00, // 247
 3.617387339134830e-01, // 248
 1.018222023184481e+01, // 249
-1.389554753911925e-04, // 250
 7.482422051278885e+00, // 251
 1.439059370704767e-06, // 252
-3.320567136524242e+03, // 253
-7.059127443743679e-02, // 254
-1.089887633368669e-02, // 255
-5.007754065873746e-04, // 256
-8.424065831272568e-03, // 257
 5.381533564797661e+02, // 258
 1.942926432299193e-03, // 259
 2.591265587215879e+01, // 260
 1.431296067963673e-03, // 261
-9.517271015586042e+00, // 262
-3.235951181676351e+02, // 263
 8.623084123084414e-03, // 264
-2.500055980982166e+02, // 265
-5.282144599454053e+01, // 266
-4.032127158068877e-02, // 267
-7.688458385087975e-01, // 268
 6.162298981061697e-04, // 269
 1.917910072106097e-04, // 270
-1.700127923674642e-01, // 271
-1.337164137118203e+02, // 272
 3.238206155651321e+01, // 273
-4.278548434802359e-04, // 274
 1.669188060518540e-02, // 275
-2.798148735023198e-03, // 276
-4.440699533578008e-01, // 277
 3.845505220131601e-04, // 278
-3.505230593140698e-07, // 279
 8.518617879243887e-03, // 280
 8.905396946978013e-02, // 281
-3.779522408107392e+02, // 282
-1.322023798677368e+01, // 283
-2.967957744254099e+02, // 284
 9.067919146690631e-03, // 285
-4.135700001347265e+02, // 286
 1.638321576467591e+00, // 287
-1.987074422079668e+02, // 288
 2.501451621513788e-02, // 289
-7.702527127044615e-07, // 290
-7.153117876409915e-07, // 291
-4.866772253258882e+02, // 292
 1.898264547092055e-05, // 293
-3.370828580335820e+03, // 294
-4.667042314701473e-01, // 295
-6.756348537200780e-01, // 296
-8.404797598657114e+00, // 297
-4.423408796128975e+00, // 298
-1.017858941626598e-01, // 299
 2.582394822661757e-04, // 300
-4.730902826744360e-01, // 301
-1.298040567116176e-06, // 302
 3.783058365777879e-04, // 303
 8.440699685426672e-01, // 304
 1.093719984200353e-06, // 305
 4.402093151378398e-11, // 306
 1.219518817052390e+03, // 307
 1.426632416172580e+02, // 308
 1.002358670357915e-05, // 309
-6.209951974303156e-03, // 310
-2.497762080981050e+00, // 311
 1.169296243025034e-04, // 312
 1.302646681631521e-05, // 313
-1.597354150619685e-03, // 314
 4.210501861609401e+00, // 315
 1.845011378662212e+03, // 316
 1.134886050624389e+01, // 317
 6.759442407974200e-03, // 318
 1.497655676027035e-03, // 319
 2.787193106270484e+03, // 320
 1.747066832106420e+00, // 321
-2.714682637299084e+01, // 322
 4.535211609339798e+00, // 323
 9.898821591030083e-01, // 324
 1.861702881984975e-09, // 325
-4.018437826836301e-03, // 326
-8.754226031527478e-04, // 327
-1.199879697352598e+01, // 328
-2.196075492190886e+03, // 329
-1.934719930460457e-02, // 330
-3.304581440135380e-03, // 331
 3.194337747077209e+03, // 332
-9.984758373614916e-01, // 333
 5.988801825079285e+01, // 334
 6.589661046816230e+00, // 335
-2.441187295511381e-01, // 336
-6.958170157133070e-04, // 337
 3.932439378844532e+01, // 338
-2.691833025290948e-08, // 339
-5.413669523811670e+00, // 340
-4.924206106116359e+02, // 341
 4.821930811136749e-01, // 342
-2.756863856481036e+02, // 343
 1.703493114724002e+03, // 344
 1.244812350583909e-03, // 345
 9.250244255910678e+01, // 346
-1.696491965538969e-01, // 347
-1.699274773212936e-01, // 348
-5.137265349659499e-03, // 349
 7.244338943001403e-01, // 350
 1.592661818453704e-01, // 351
 4.313324036932629e-01, // 352
 3.602861278961067e-04, // 353
-2.611109335838023e-01, // 354
 5.070639763092572e+00, // 355
 7.632638375341045e-03, // 356
-7.673981934556191e+01, // 357
 4.934959855265739e-01, // 358
 9.248281067734657e-05, // 359
 3.900168964026963e-06, // 360
-1.504394521728031e+02, // 361
-1.412173872644945e-01, // 362
-6.172283826057150e-11, // 363
 6.119944054504032e-01, // 364
 1.091044619894167e+03, // 365
-3.654157375418982e+02, // 366
 1.370607090781435e+00, // 367
-1.351311003545443e+03, // 368
 2.542449040549704e+03, // 369
-1.295581149979607e-06, // 370
 8.376274423767806e+01, // 371
-3.271657989037155e-01, // 372
 2.108104827992628e-01, // 373
-7.925685162854832e-03, // 374
-2.903958868402133e-06, // 375
 1.910194001389095e+03, // 376
 1.075658314255070e+03, // 377
 1.297551613944612e+03, // 378
 1.758942327097579e+02, // 379
-2.252525563289825e+03, // 380
-9.813422796840159e-01, // 381
-6.643318897295769e-01, // 382
-7.691368614758642e-01, // 383
-1.445584757875615e-02, // 384
 5.055988266739043e+02, // 385
-7.592696256932015e+02, // 386
-2.627455087911121e-01, // 387
 2.527934691705224e-02, // 388
-6.452853915763633e+02, // 389
 1.994389793762115e+02, // 390
 1.141893501458339e-04, // 391
-1.122396052656554e-06, // 392
 5.637718993978204e-10, // 393
 1.348972198304682e-04, // 394
-3.040993462953917e-04, // 395
-1.491533406605193e-04, // 396
 1.248614631123028e-02, // 397
-4.725943216171859e-02, // 398
-3.472444821620171e+01, // 399
 4.089307174747211e-06, // 400
 6.948897866893716e-01, // 401
-5.153795468315222e-01, // 402
 7.758366434243013e+01, // 403
-2.717503397288142e+00, // 404
 1.177691299048881e-06, // 405
 4.992732693947232e-02, // 406
 5.604008066831983e-03, // 407
-3.134904815298161e-04, // 408
 1.399147942566751e+01, // 409
-1.195435489256700e-03, // 410
 1.603096578837707e-06, // 411
 1.614143682110456e+01, // 412
 1.974487553626041e+00, // 413
 4.687558316137558e+02, // 414
-8.015342168505667e-02, // 415
 1.346109939160783e-01, // 416
 2.222732746835571e-02, // 417
 1.240128565692754e+02, // 418
-1.244936102222522e-04, // 419
-8.946658684911072e-03, // 420
-5.227310602310110e-01, // 421
-1.032292495616846e-07, // 422
-2.093054691297406e-02, // 423
-3.429377247806899e-09, // 424
 3.822106519234097e+02, // 425
 4.152575754600822e+02, // 426
 1.044192172182904e-08, // 427
-3.922067753875728e-02, // 428
-2.270704146918421e-02, // 429
 2.693873237432851e+01, // 430
 3.521378669993908e+00, // 431
-4.782705392250661e+01, // 432
 3.144494538280628e+02, // 433
 1.338170303218184e-06, // 434
 6.717480112285018e-02, // 435
 7.302898073005912e-01, // 436
-4.158830059186869e+02, // 437
 5.361571245563300e-03, // 438
 6.056921039780614e+02, // 439
 5.331412253967022e-01, // 440
-2.939254361419780e-01, // 441
 9.265719184823355e+02, // 442
 3.932256296477937e+01, // 443
 1.916941518260488e-04, // 444
-1.174783425843209e-02, // 445
-1.883302734502256e+02, // 446
-5.954934601975332e-02, // 447
 9.104411402458492e-03, // 448
 2.191725011326147e-01, // 449
-1.565702155022452e+03, // 450
 1.822367227176060e+01, // 451
 7.051519360064599e+00, // 452
 1.141442928490812e+01, // 453
 1.604265415758033e+00, // 454
 8.329769511844926e+02, // 455
-9.630325842287514e-03, // 456
 7.006138540560472e+02, // 457
 2.837889172345702e-04, // 458
-2.107473358977351e-01, // 459
 1.463129592987357e+03, // 460
 7.839753866218440e+02, // 461
 6.065557365621867e+02, // 462
 3.280958113925359e+01, // 463
 8.954304243459841e+02, // 464
 4.824345016111154e+02, // 465
-4.767986696906407e+02, // 466
 5.609753101223049e-01, // 467
-1.425081107418690e+01, // 468
-4.571642633697629e-05, // 469
 3.051751696700950e-09, // 470
-2.544900860336775e+00, // 471
-5.015969182743870e+01, // 472
 1.374496395642898e-02, // 473
 1.430447401466606e-02, // 474
 4.031503490837629e+02, // 475
 1.015015187937611e+01, // 476
 4.638514760103257e-05, // 477
 1.622136784557067e+02, // 478
 9.848686805517113e+01, // 479
 2.303628287893098e+00, // 480
-2.440017829307484e+03, // 481
 2.353561947305212e+03, // 482
 1.154416383023976e+03, // 483
 3.371253403430238e+02, // 484
 4.077980584387028e+03, // 485
-1.189520919770826e-04, // 486
 3.141729444994834e+02, // 487
 5.280839919075211e+02, // 488
-1.012058475652642e+03, // 489
 7.307784876214833e+00, // 490
 2.670683388973212e+03; // 491

}
