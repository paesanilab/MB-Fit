netcdf x2b_A1B2_A1B2_v1x {
  // global attributes 
  :name = "x2b_A1B2_A1B2_v1x<4>";
  :d_intra_AB =  2.983850399822167e+00; // A^(-1))
  :k_intra_AB =  1.999779699119901e+00; // A^(-1))
  :d_intra_BB =  2.765428437998016e+00; // A^(-1))
  :k_intra_BB =  1.999999644482479e+00; // A^(-1))
  :d_AA =  2.434958510788339e+00; // A^(-1))
  :k_AA =  2.615539497340414e-01; // A^(-1))
  :d_AB =  4.276801423395641e+00; // A^(-1))
  :k_AB =  1.351515115768721e+00; // A^(-1))
  :d_BB =  4.148041188197417e+00; // A^(-1))
  :k_BB =  1.770346740483469e+00; // A^(-1))
  :r2i =  6.000000000000000e+00; // A
  :r2f =  7.000000000000000e+00; // A
  dimensions:
  poly = 597;
  variables:
    double poly(poly);
data:
poly =
-1.716556897235306e+02, // 0
 1.879151260546268e+02, // 1
 5.039820869809339e+02, // 2
-1.247827758917015e+02, // 3
-3.866091164586685e+01, // 4
-1.297231571887610e+01, // 5
 6.511917877329410e+00, // 6
 1.834097571700555e+02, // 7
 1.201999652181833e+01, // 8
 1.155959329946990e+02, // 9
-2.162259508967571e+00, // 10
-4.886238825430601e+00, // 11
-1.563406968957204e+01, // 12
 1.238154368960775e-01, // 13
 1.414111524612345e+00, // 14
 5.162978113410981e+01, // 15
 1.719733640880105e+00, // 16
 7.003010529204444e+00, // 17
-2.402082549429714e+00, // 18
-2.252918284504474e+00, // 19
 2.157367480830090e+02, // 20
-2.254059332791383e+00, // 21
 6.829252268675213e-01, // 22
-4.652994917947478e+02, // 23
 9.300558520711808e+00, // 24
-8.138593481886010e-02, // 25
-5.792019186792743e-04, // 26
 7.786071618844005e-02, // 27
-3.916143432353687e-03, // 28
-1.610474914152116e+00, // 29
 1.777978318982538e-01, // 30
-3.439263946981387e+00, // 31
-3.741438268105712e-02, // 32
 1.387228489850003e-01, // 33
 2.094031362571654e-02, // 34
-3.154917292036287e+00, // 35
-3.154713773299916e-02, // 36
 1.994322638997634e-02, // 37
-2.186413294865106e-01, // 38
 4.168126579199391e+00, // 39
 1.964113168248353e+00, // 40
 4.230081395329690e+01, // 41
 7.561233555780326e-02, // 42
-2.467953085365694e+00, // 43
 4.726662856919633e+00, // 44
 8.620594623710136e+01, // 45
 2.031928855070474e-02, // 46
-2.448659914796902e-01, // 47
-1.508949689825486e+00, // 48
-2.412848641816323e+00, // 49
-4.213323037050877e-04, // 50
-1.925236767338710e-04, // 51
 2.294596219566061e-01, // 52
 8.078133630818069e-03, // 53
-4.116006054938521e-03, // 54
-1.070048223672037e-01, // 55
-1.366547524102005e+01, // 56
 7.704753234564004e-01, // 57
 9.670851979328873e-01, // 58
-1.027357006069268e-02, // 59
-3.341990969833170e-03, // 60
 3.032849493363427e+02, // 61
-4.413447971460323e-02, // 62
 1.976873511964267e-01, // 63
 2.422295682093698e+00, // 64
 2.703440729320113e-02, // 65
 2.361129284689498e+01, // 66
 7.374646694548200e-03, // 67
-1.010284354453870e+01, // 68
-1.212972753576132e-02, // 69
-1.724225384884444e-01, // 70
 2.813195642610650e+00, // 71
-2.786654700579660e+00, // 72
-1.816703782794628e-01, // 73
-1.141103025305116e-02, // 74
-1.499695761831053e-01, // 75
 8.041844007803198e-02, // 76
-2.818473816781513e-02, // 77
 1.640408108926979e-02, // 78
-1.097444456972649e-01, // 79
-2.455372265214589e+01, // 80
 2.989571981305021e+00, // 81
-1.282312783787553e-01, // 82
-1.887195329536906e-02, // 83
-5.378502966956154e-04, // 84
 2.069239571007967e+01, // 85
 7.375050683753599e-02, // 86
 6.064473925663631e+00, // 87
-2.930977583604875e+01, // 88
 4.044037472940169e-01, // 89
-3.093884103164986e+00, // 90
-7.467497673243489e-04, // 91
-3.754036318309316e+00, // 92
-2.636940124269609e-03, // 93
-1.396212489603397e+02, // 94
-1.794071829628349e-03, // 95
-4.485740334338928e-02, // 96
 2.579452398815667e-02, // 97
 9.543199100665294e-02, // 98
 1.481164407861118e-01, // 99
-6.372825337270904e+00, // 100
 2.469403412423648e+00, // 101
-4.252842387855442e-03, // 102
-7.549207034841650e-02, // 103
-1.688579849190709e+01, // 104
 4.814117795205982e-01, // 105
-2.556409534402539e+00, // 106
-1.203728613974232e+00, // 107
 5.763846810508688e-01, // 108
-3.450186694201782e-05, // 109
 2.179550133610488e+01, // 110
-2.660242955459958e-03, // 111
 7.281028453722113e+00, // 112
-2.152150134279503e+01, // 113
 9.270142955439552e-02, // 114
-8.269122120858768e-02, // 115
 2.594620240835611e+00, // 116
 7.110361026248326e+01, // 117
 1.128092640861917e-01, // 118
 1.674763206907787e-01, // 119
 7.165602112330489e-02, // 120
-4.580988280904382e+00, // 121
 3.940267891972088e-03, // 122
-9.925981076187562e-02, // 123
 9.289465048767491e-01, // 124
-8.243869262619506e-02, // 125
-3.208296887230917e+01, // 126
 3.059615457414176e+01, // 127
-3.493249444708971e+00, // 128
-5.793668015057370e+00, // 129
-1.396305205607103e+01, // 130
-9.218144313130595e-03, // 131
 8.659201071758957e-01, // 132
-1.097819825925450e+02, // 133
-6.845367056058764e-05, // 134
-2.340635706608816e-01, // 135
 3.167087989016046e-02, // 136
 1.686669226980191e-04, // 137
-5.214077148121619e-02, // 138
 3.185177936333270e-05, // 139
 9.453893369733830e-05, // 140
 1.360097341380329e-04, // 141
-2.461013286042055e-01, // 142
-1.908709733590772e-03, // 143
 1.600419597162766e-03, // 144
-9.861074842552597e-08, // 145
 1.707020549020515e+00, // 146
 1.434892774487877e-03, // 147
 5.867310950075670e-04, // 148
 8.931414649290836e-05, // 149
 2.793693789577585e-01, // 150
-5.894243284284279e-04, // 151
 1.722341753915645e-04, // 152
-1.684894745386747e-02, // 153
-2.808810718777621e-04, // 154
-1.057143256133141e-04, // 155
 5.920317342252019e-04, // 156
-6.325496558657866e-05, // 157
-1.426166430586631e-02, // 158
-1.214727109215763e+00, // 159
 2.599183561161458e-05, // 160
-9.600336266323516e-03, // 161
-3.835600415125575e-02, // 162
-1.236599678920506e-03, // 163
 4.493970700629176e-03, // 164
 5.235990430156014e-03, // 165
-2.918898540694079e-01, // 166
-7.015079673282481e-04, // 167
 5.692873354994837e-02, // 168
-2.363060211678033e-06, // 169
 1.605740391675895e-03, // 170
-3.989126306642274e-04, // 171
 1.272253698587554e-01, // 172
-2.957782142076314e-02, // 173
 3.354171128806122e-01, // 174
-1.226385053387462e-03, // 175
 1.653980811824546e-04, // 176
 1.874899497428916e-02, // 177
 9.524671818597293e-04, // 178
 4.569022482840719e-02, // 179
-8.707477877345283e-04, // 180
-1.832903706476481e-04, // 181
 9.029080984329462e-03, // 182
-2.112892089252288e-01, // 183
-2.797362238459848e-02, // 184
 3.068172650321364e+00, // 185
 4.936938992109156e-05, // 186
 1.613366889360247e-03, // 187
-9.219338728173769e-05, // 188
 7.480388382199693e-05, // 189
 3.530811327947373e-02, // 190
-5.800254416857796e-03, // 191
 2.796363359004159e-03, // 192
-9.942654172732066e-05, // 193
-2.925607541472559e-01, // 194
 1.958670105927303e-05, // 195
-7.271329659492531e-04, // 196
-1.839449611990414e-04, // 197
-3.533493681076704e-01, // 198
 1.418185634663058e-05, // 199
-7.540633031241515e-05, // 200
 8.694590947126456e-05, // 201
 1.490048998589548e-05, // 202
 2.968094047701594e-02, // 203
-1.850277404876925e-05, // 204
 5.911221573551778e+00, // 205
-5.164990782462965e-06, // 206
 4.832370891541226e-05, // 207
-7.561384824525854e-04, // 208
 2.705930176162145e-01, // 209
-3.063491556071393e-06, // 210
-2.206762251433561e-02, // 211
-1.337856521981954e-01, // 212
 4.907056265338213e-05, // 213
 2.333094169204108e-05, // 214
-9.858314226182447e-01, // 215
-1.435317466762683e-04, // 216
-2.584107629693371e+00, // 217
 2.096324391450464e-02, // 218
 8.248082435330717e-02, // 219
-1.669036232234631e-03, // 220
-1.855619534960070e+00, // 221
-2.570027972477456e-05, // 222
 2.444783095784150e-02, // 223
-1.742275677487474e-06, // 224
 2.459018064955142e-02, // 225
-1.278228400862733e+01, // 226
 1.331518323338379e-01, // 227
-2.564792621944090e-03, // 228
 1.738127782446646e-05, // 229
-7.557151013433652e-03, // 230
-2.717710313579807e-06, // 231
 3.654629356064382e-03, // 232
 7.836173440672303e-06, // 233
-3.166458428978239e-06, // 234
-1.397378050605858e-03, // 235
 2.892807435598958e-06, // 236
-7.544842248782194e-02, // 237
 9.560580528319643e-01, // 238
-1.421032696137721e-06, // 239
-3.595892077194916e-07, // 240
-3.587091941078395e-02, // 241
-1.575210778934655e-01, // 242
 1.589495143204839e-03, // 243
-1.083383591842908e-04, // 244
 3.388767958482669e-01, // 245
-4.737433716126536e-05, // 246
 1.442261876850306e-03, // 247
-2.962775526169499e-03, // 248
-2.371003560192524e-03, // 249
-6.080167467079466e-05, // 250
 1.368822131962558e-02, // 251
 4.180225375746448e-06, // 252
 5.157717145380287e-05, // 253
 1.818285965041310e-06, // 254
-5.526941693902825e-06, // 255
-2.425862093088478e+01, // 256
-1.199555859068424e+00, // 257
 6.977111473707100e-01, // 258
-1.864028892068867e-04, // 259
 2.007286274561204e-01, // 260
-4.288902746732647e-04, // 261
-9.298757516551258e-04, // 262
 8.272056090804499e-03, // 263
 9.481927027465004e-03, // 264
-2.775210943656346e-02, // 265
-1.607812280127022e+00, // 266
-9.190836056382041e-05, // 267
-6.430908344326504e-03, // 268
-1.052151831320898e-03, // 269
 7.113331005877642e-05, // 270
-9.799055436629121e-02, // 271
-5.227855244124453e-04, // 272
 8.393855620257416e-07, // 273
-3.138605763056356e-01, // 274
 2.126626350286886e-03, // 275
 1.032951595035188e-03, // 276
 9.381768613643589e-03, // 277
-1.545283067935578e-01, // 278
-7.567043754144994e+01, // 279
 1.361763333062771e-02, // 280
 8.408143512519385e-06, // 281
 3.973326370029298e-04, // 282
 8.295562759508307e-02, // 283
 9.156916153046516e-01, // 284
 4.591406898801763e-03, // 285
-1.429589996222311e-04, // 286
 2.171213553741199e-02, // 287
 1.677686926815961e+01, // 288
 5.682693930254928e-02, // 289
-7.591560306332474e-01, // 290
-2.213253185838960e-06, // 291
-4.354608201197662e-03, // 292
-1.567387484161371e-01, // 293
 4.784118395112894e-05, // 294
-9.479932126827663e-02, // 295
-1.741649847104552e-02, // 296
 3.006376791456373e-02, // 297
-1.735945141469909e-02, // 298
 2.779525440484528e-08, // 299
 1.930372336074253e-02, // 300
-3.185896627122045e+00, // 301
-3.438530575888692e-01, // 302
-1.293400780967018e-02, // 303
-3.442203636828777e+01, // 304
-3.370419646142632e-04, // 305
 2.919745502010507e-03, // 306
 2.158956557511066e-06, // 307
 1.306190441304346e-03, // 308
-1.555306291334068e-02, // 309
 1.890336838631501e-04, // 310
-2.576747704932937e-03, // 311
 1.369012638218179e-01, // 312
 4.778181188099120e-02, // 313
 2.650027875984412e-05, // 314
 4.411340154513270e-03, // 315
-4.105357431822321e-06, // 316
 1.070426846355015e-03, // 317
 9.707381478897539e-03, // 318
 1.068583201964382e-03, // 319
-3.361311983835621e-03, // 320
-8.217635257488888e-02, // 321
 2.475549838594093e-03, // 322
 4.979672205429569e-02, // 323
 2.581196611328174e-05, // 324
-1.220649672675155e-05, // 325
-1.690393042377430e-04, // 326
 3.384329176766537e-01, // 327
 3.746192708830797e-02, // 328
 6.902909962174275e-02, // 329
-1.071529407998110e-03, // 330
 2.858365230584651e-03, // 331
 2.562017688877905e-04, // 332
 1.352841028831073e-04, // 333
-9.881533769351825e-01, // 334
-8.653232237567658e-01, // 335
-6.974304374693823e-03, // 336
-3.986532618007387e-01, // 337
 3.012844167148236e-05, // 338
-6.716315923557909e-05, // 339
 2.446699086243252e-02, // 340
-8.233849812945032e-04, // 341
 6.458384908023714e-02, // 342
 1.001751049671995e-01, // 343
 9.573634891336282e-04, // 344
-4.312771427229777e-04, // 345
-3.957248616381775e-04, // 346
-5.874678835477386e-02, // 347
 4.600823735596485e-01, // 348
 2.203908586096169e-06, // 349
 7.113477060778529e-03, // 350
-6.396974921586585e-02, // 351
 1.342579781042404e-01, // 352
 1.074355660789059e+01, // 353
-8.091359805978551e-03, // 354
-4.808228389771373e-02, // 355
 5.754394449492544e-02, // 356
 1.419396519221854e-05, // 357
-3.175463427718980e-02, // 358
 2.325812327953980e-02, // 359
 1.399833964563963e-01, // 360
-1.134368810404512e-01, // 361
 7.671215286322756e-02, // 362
 1.466733697778382e-03, // 363
 2.078212448892627e-05, // 364
 4.458984479165855e-06, // 365
-1.362919790981182e-02, // 366
-4.083337722194927e-05, // 367
-1.074470167306995e-04, // 368
-2.132109010305891e-02, // 369
-4.906484777805555e-03, // 370
 9.816315723924289e-03, // 371
-9.620024744633882e-07, // 372
 1.040329271867847e+00, // 373
-1.968914728616670e-04, // 374
 1.273562953541104e+00, // 375
-9.157843664723067e-02, // 376
-6.357108824302319e-05, // 377
-9.324268977176340e-06, // 378
-4.316421164855571e-05, // 379
 8.241741814985059e-03, // 380
 5.060593751900285e-03, // 381
-7.804380568685685e-04, // 382
-1.065223542622957e-02, // 383
-2.745890878405603e-02, // 384
-2.320052897183116e-03, // 385
 2.964231586246738e-04, // 386
-2.327207344992142e-03, // 387
-2.039260578648690e-05, // 388
-8.791021380004012e-07, // 389
 1.898672664124969e-04, // 390
 1.327228839198776e-05, // 391
-1.770654998637529e-02, // 392
-1.974407468415484e-06, // 393
-1.509407810344513e-05, // 394
 3.165982675073240e-03, // 395
-1.387944689065637e-04, // 396
-9.242126242332525e-05, // 397
 8.360299825364483e+01, // 398
 1.208640046412657e-03, // 399
-1.085384425503120e-03, // 400
 5.840433416499413e-04, // 401
 3.059113364152188e-01, // 402
 5.145873886430700e-05, // 403
 1.008019653951814e+00, // 404
 1.113116874963745e-02, // 405
 2.240862594544266e-03, // 406
-8.337597661717002e-01, // 407
-1.616395854567543e-03, // 408
-1.442956856550336e-02, // 409
 5.612066166425459e+00, // 410
-1.726278252972622e-04, // 411
 7.675776402387301e-06, // 412
-6.736876003965535e+00, // 413
-1.297178158508013e-02, // 414
 1.970897378224283e-03, // 415
 3.526372191139374e-02, // 416
 3.791888016222354e-02, // 417
-1.068306741693274e-02, // 418
 1.580693932292379e-03, // 419
 1.041984688085287e-03, // 420
 1.036350639803806e-04, // 421
 4.617065922110100e-06, // 422
 2.227736763922636e-02, // 423
 8.262406667217208e-04, // 424
 1.296557522813072e-03, // 425
-1.213100034499293e-04, // 426
-4.558869953765917e-02, // 427
 1.011614966043334e-05, // 428
 4.943008423531791e-05, // 429
-1.623232010991195e-02, // 430
-9.289874531234971e-05, // 431
-1.511531820257878e-06, // 432
-5.050550758799437e-04, // 433
 3.689390687584710e-02, // 434
 1.745531495652201e-04, // 435
 2.435716518136707e-06, // 436
 2.076218603511612e-06, // 437
 7.723680001748195e-01, // 438
 1.046606919584248e-03, // 439
-3.036422777092234e-02, // 440
-3.740787986820641e-02, // 441
-6.610876927255221e-05, // 442
 4.557037058104172e-03, // 443
 3.722276651069834e+00, // 444
-6.416008658678002e-05, // 445
-6.397845306130731e-01, // 446
-4.804911980766702e-03, // 447
-8.639482190739733e-04, // 448
-6.297967754380288e-05, // 449
 8.348954928128662e-05, // 450
-6.920351203643164e-01, // 451
-3.153605003385474e-05, // 452
 3.581200363239791e-03, // 453
-9.838515213635657e-01, // 454
 1.182414318179773e-06, // 455
-9.059518566003353e-03, // 456
 1.866695154604298e-02, // 457
 1.957538624139961e-03, // 458
-6.424799195826356e-06, // 459
-2.588387371005352e-03, // 460
-1.444425707368094e-01, // 461
-5.247427458823497e+00, // 462
 3.504363377532827e-04, // 463
-6.413250131101013e-04, // 464
 1.949970412096430e-03, // 465
-1.323207212693686e-01, // 466
 8.716499271409281e-01, // 467
-9.961408991564033e-05, // 468
 1.456615747864683e-01, // 469
 3.378280013983919e-03, // 470
 1.777600687530090e+00, // 471
-1.900942511757328e-03, // 472
-4.646922485074021e+00, // 473
-8.656952812762039e-04, // 474
-1.999100895000587e+00, // 475
-5.502560675973222e-04, // 476
-9.615162959959268e-06, // 477
-3.444363999407403e-03, // 478
 1.312038210004132e-03, // 479
-6.280301018567329e-06, // 480
 1.140833537843744e+01, // 481
 1.711707128581770e-06, // 482
-2.319982453842070e-03, // 483
 2.431914025291860e-03, // 484
 3.153426569902579e-02, // 485
 9.532190376515748e-05, // 486
-9.038622693494143e-06, // 487
-3.640765294624636e-02, // 488
-9.092811005227076e-02, // 489
 1.236002012935657e-05, // 490
 8.103495734631592e-01, // 491
 2.207072643150293e+01, // 492
 1.422367755041600e-04, // 493
 8.523306171444551e+00, // 494
 1.142081307736496e+00, // 495
-1.407280969489307e-04, // 496
 3.036382402139211e-05, // 497
 3.291131205653565e-02, // 498
 1.295327623846089e-01, // 499
-6.376102262590329e-02, // 500
-6.113916619403766e-04, // 501
-8.916784036483258e-06, // 502
-4.485142629465583e-06, // 503
 1.996345271836891e+00, // 504
 1.129636277927699e-05, // 505
-1.473110843263368e-04, // 506
 1.486111802277672e+00, // 507
-1.922241630532361e-07, // 508
 9.862100381488883e-04, // 509
 2.692674838450866e-04, // 510
 2.414537270534907e-04, // 511
 4.514253844873805e-05, // 512
 8.940004757937716e-03, // 513
 2.572771072267381e-02, // 514
-6.092337581904431e+00, // 515
 5.290540224845828e-06, // 516
 1.043763609017330e-06, // 517
 9.488746135755683e-06, // 518
 2.828347327551668e-05, // 519
 1.129464769528758e-04, // 520
-1.330687050976488e-04, // 521
-9.717669667554876e-02, // 522
 1.685814886599643e+00, // 523
 9.099582157861275e+01, // 524
 3.326833551968641e-05, // 525
 2.230705762425298e-03, // 526
 2.053523960172086e+01, // 527
 3.196261964409918e-01, // 528
 8.186826151278916e-01, // 529
 2.787258937880249e-04, // 530
 1.066760503721308e-01, // 531
-3.227629489922871e-01, // 532
 7.857085391641105e-03, // 533
-2.237646025739057e+01, // 534
-8.591588253781215e-03, // 535
-1.169229553700476e-03, // 536
 1.067840227833299e-01, // 537
 4.937406768025969e-01, // 538
 9.658059945917240e-04, // 539
 1.302086066023000e-04, // 540
-3.415639682760944e-02, // 541
-1.024820422084977e-04, // 542
-1.750694353049260e-06, // 543
 4.979303690931365e+00, // 544
-1.623631515250796e-04, // 545
-4.398202359113392e-06, // 546
 2.292847386483875e-03, // 547
 2.978469014827690e-04, // 548
-1.536156175551862e+00, // 549
-3.216623651819265e-06, // 550
-3.548299972482152e-05, // 551
 3.497867377058236e-02, // 552
 8.932108589243422e+00, // 553
 3.004801963780915e-02, // 554
 4.681206556502806e-03, // 555
-7.231452219408710e+00, // 556
 2.542990212624920e-02, // 557
-2.066348012677322e+00, // 558
 8.170163805235046e-04, // 559
-1.171408137317913e-03, // 560
-1.387351787694429e-03, // 561
-8.106323493577346e-02, // 562
-2.642228287830767e-03, // 563
 9.314685409035576e-03, // 564
-6.423008286943603e-04, // 565
 1.121321652476487e-05, // 566
-3.774204697288546e-03, // 567
-3.897751724105811e-02, // 568
 4.251127412567280e-02, // 569
-4.023485684598991e-01, // 570
 4.940717430351327e-05, // 571
 1.408520841752720e-03, // 572
 6.189189464693792e-02, // 573
-1.366335960653411e+00, // 574
 1.053356164165175e-05, // 575
 1.856942045638767e-06, // 576
 1.547761521667615e-02, // 577
 6.514090081965193e-05, // 578
-8.177835088265077e-02, // 579
 1.827959599135587e+00, // 580
 2.170631199402664e+00, // 581
 2.320327730432315e-01, // 582
-5.382135566064016e-01, // 583
-2.965185704952006e-06, // 584
-2.741732314115159e-03, // 585
-1.628387972842725e+00, // 586
 2.396104807804857e-05, // 587
-1.069076487850218e-03, // 588
-1.420233493118088e+02, // 589
 1.365104506088591e+00, // 590
 1.818438862020880e-02, // 591
-7.259791180535294e-02, // 592
-4.587868589411698e-03, // 593
-1.556950079770190e-04, // 594
 1.832091173177896e-01, // 595
-2.522450271681962e+02; // 596

}
