netcdf x2b_A1B2_A1B2_v1x {
  // global attributes 
  :name = "x2b_A1B2_A1B2_v1x<4>";
  :d_intra_AB =  3.078705151200680e-01; // A^(-1))
  :k_intra_AB =  5.711075064676757e-01; // A^(-1))
  :d_intra_BB =  2.598399713421982e+00; // A^(-1))
  :k_intra_BB =  3.914551121181958e-01; // A^(-1))
  :d_AA =  1.062122784836762e+00; // A^(-1))
  :k_AA =  2.992028280624167e+00; // A^(-1))
  :d_AB =  1.544504632076253e+00; // A^(-1))
  :k_AB =  3.898082729747417e-01; // A^(-1))
  :d_BB =  3.171873714136767e+00; // A^(-1))
  :k_BB =  2.996623286333546e+00; // A^(-1))
  :r2i =  6.000000000000000e+00; // A
  :r2f =  7.000000000000000e+00; // A
  dimensions:
  poly = 597;
  variables:
    double poly(poly);
data:
poly =
 2.550638499287735e+02, // 0
-2.496008640769404e+02, // 1
 6.706357378617221e+02, // 2
-5.133983206333849e+02, // 3
 2.085350421967280e+02, // 4
 5.408028940892591e+03, // 5
-1.523906275218335e+02, // 6
-3.909774644334291e+03, // 7
 6.611915658837653e+03, // 8
-6.632315536041468e+02, // 9
 3.890073273855485e+02, // 10
-1.478709203290974e+02, // 11
 3.154710965074879e+00, // 12
-1.440406466497513e+00, // 13
-6.696684914900988e+03, // 14
-2.244026532766819e-01, // 15
 1.815308680941738e+01, // 16
-4.863621613170223e+03, // 17
 4.469325209611165e+03, // 18
 1.835333351296725e-01, // 19
 4.560174547392106e+02, // 20
-4.317345841190575e+03, // 21
-2.121287646568573e-01, // 22
 1.428213336641075e+04, // 23
 3.196263328381483e+02, // 24
-3.684784741476538e+03, // 25
 2.580251496353903e-04, // 26
 5.243183355154108e-01, // 27
 5.002562012666191e-01, // 28
 2.296901511719444e+01, // 29
 3.766964347316311e+02, // 30
 1.786993772771295e+03, // 31
-1.355100104592890e+00, // 32
-6.150096995162407e+03, // 33
 1.479788626527779e+01, // 34
 1.621911795833115e-01, // 35
-7.804546564923077e-03, // 36
 1.921386599165860e-01, // 37
-5.393884005753181e+01, // 38
-2.357676254324267e+03, // 39
-3.300827660536750e+03, // 40
 5.931477610914608e+03, // 41
 5.398263137267403e+02, // 42
 1.218479467889711e+00, // 43
 1.060706741189181e+01, // 44
-2.374641384996211e+03, // 45
 4.103145294786866e+01, // 46
 8.635717854538291e+02, // 47
-2.412523782196835e+00, // 48
 3.156276377702514e+01, // 49
-3.494236499571453e-05, // 50
-5.101716667373113e+03, // 51
 7.015369435542816e-01, // 52
-1.360061088244272e+01, // 53
 2.060232112433114e+00, // 54
-5.494935662786937e+03, // 55
-3.817680851483329e+02, // 56
-3.075483529526417e-01, // 57
 2.951455539773007e+00, // 58
-2.236133790686047e-03, // 59
 8.261264905645698e+03, // 60
-3.594975909105153e+01, // 61
 7.608545366918873e+03, // 62
-5.960512117395971e+01, // 63
 4.435410261778799e+03, // 64
 1.355564676947680e+01, // 65
 8.146764001789831e-01, // 66
 4.142960854756104e-01, // 67
-2.168589377349332e+02, // 68
-4.150458108570763e+03, // 69
-1.101347116544747e+01, // 70
 4.004911887517346e+03, // 71
 1.569530647658466e+03, // 72
-2.416729351031933e-02, // 73
 5.397004727137090e+03, // 74
-1.515174750663035e+02, // 75
-2.406821396277920e+02, // 76
-2.882785073865274e+01, // 77
-2.950294960391266e+00, // 78
-1.377331512302197e-03, // 79
-3.638912163474059e+01, // 80
 4.065728952127790e+03, // 81
-8.358908392126042e-02, // 82
 2.176930404358118e+00, // 83
-1.158773837142620e-03, // 84
-2.494474139241885e+03, // 85
-4.401203791334574e+03, // 86
-1.244395072090470e+02, // 87
-5.437539248733445e+02, // 88
-8.095848939076821e+01, // 89
-5.795695391157190e+03, // 90
 6.283834442835857e-03, // 91
 8.327287430612784e+02, // 92
-4.139364542960524e+03, // 93
-1.014518819714597e+03, // 94
-1.344337005111068e+01, // 95
 3.556973423718626e+03, // 96
-1.387073193452503e+01, // 97
 3.695943545153984e+02, // 98
 1.705828661362185e+01, // 99
-3.124125140956008e+03, // 100
-6.880344696281903e+03, // 101
 2.691679711034104e+02, // 102
-1.693202333892439e+02, // 103
-5.584210867974464e-06, // 104
-2.903495816935003e+02, // 105
-5.316877090121697e+03, // 106
 1.127361465781776e+04, // 107
-2.624851875749782e-04, // 108
 2.255366544420498e+00, // 109
 3.834341642595431e+02, // 110
 8.017179386196512e+03, // 111
-1.269709640030514e+03, // 112
-3.738233350726905e-01, // 113
-1.695431348198130e+04, // 114
 2.627433212130741e+00, // 115
-5.775710319683379e+02, // 116
-2.810408725112005e+01, // 117
-2.154857918207440e-04, // 118
 3.034323645754981e+03, // 119
 5.179999038042245e+03, // 120
 1.052311864455351e+04, // 121
 9.756597941527810e-02, // 122
 3.352528449611440e-06, // 123
-7.235253190402936e+03, // 124
-1.102609930336223e+03, // 125
-2.103713178725343e-02, // 126
 3.894804023133048e+03, // 127
 2.416261362808126e+03, // 128
 2.988381910749606e+00, // 129
-1.584551208199793e-02, // 130
-3.376009379976696e+02, // 131
-5.930339921383387e-01, // 132
-3.411497638865302e+03, // 133
-6.987556656641916e-02, // 134
 1.003380204193312e+03, // 135
 1.961742260191193e-01, // 136
-1.160264236943521e-04, // 137
 2.815392836650689e+00, // 138
-7.319831898620484e-04, // 139
 1.704193614713486e-03, // 140
 2.750639688896170e+01, // 141
 3.927023750948722e+03, // 142
-6.002420205884119e+00, // 143
 5.466141951080728e+01, // 144
-3.110966268651522e+00, // 145
 6.742054158190036e+02, // 146
-4.920287636799484e-03, // 147
-2.966765775283601e+01, // 148
 1.288905017162551e+00, // 149
-1.437434662712287e+02, // 150
-2.188780776166522e-04, // 151
-6.238847748764866e-01, // 152
-1.255844200504439e+03, // 153
-4.247718563648794e-01, // 154
-3.429825405888506e+01, // 155
-5.802287087118599e-04, // 156
-4.148538907881538e-01, // 157
 1.345745814796768e+01, // 158
-2.521792692989073e+03, // 159
 2.130437944451127e-04, // 160
-1.019498054623961e+02, // 161
-3.347683399528633e+00, // 162
 2.124314672461566e-03, // 163
 5.440819204345137e+01, // 164
 8.703302362825418e+02, // 165
-8.968278811336989e-01, // 166
 1.742088744871587e-03, // 167
-3.876348658791503e+03, // 168
-1.424004293634606e-06, // 169
 4.111939269563262e+03, // 170
 9.843965620262925e-04, // 171
 5.056144879910264e+01, // 172
 5.137991015232210e+03, // 173
 9.560260464373971e+03, // 174
-8.832980297135895e-04, // 175
-5.349278237433894e-03, // 176
 1.534722663478778e-01, // 177
 3.321281672594177e+03, // 178
-5.820847287642374e+00, // 179
 1.911397393173524e+03, // 180
-3.068138822192763e+01, // 181
-8.069168936167977e+02, // 182
-4.361270558389089e+01, // 183
-6.932388713064914e-02, // 184
-1.279705747427823e+00, // 185
 1.613025957450219e+03, // 186
 2.145712319939229e-02, // 187
 5.576907696082621e-04, // 188
-1.255656018098841e+00, // 189
-2.811300331520771e+03, // 190
-9.697704548868121e-01, // 191
-9.211189493901732e+01, // 192
 1.093950167775574e+01, // 193
-1.937553506378215e-05, // 194
 3.265293496708252e+01, // 195
-4.073740138615664e+03, // 196
 1.515282746132376e-04, // 197
 1.804961804298186e+00, // 198
 3.776422806701303e+03, // 199
 4.822853543915648e-02, // 200
-2.068330586794627e-06, // 201
-2.397189657289714e+01, // 202
 2.126981947652300e+00, // 203
-1.399363429668450e+02, // 204
-7.711376990403702e+02, // 205
 7.590162217929393e-01, // 206
 6.954864330202185e-07, // 207
-6.163250055067745e+03, // 208
 2.254697836505830e+00, // 209
 3.485593339935241e+00, // 210
-1.632065054822941e-02, // 211
-6.836489665860586e-02, // 212
-4.703911476436953e+03, // 213
-3.136345824953719e+00, // 214
-1.423128593054149e+01, // 215
 1.134246489818477e+00, // 216
-9.423363357890164e+00, // 217
 8.420830260625696e+00, // 218
 9.062308220588650e+02, // 219
-7.899555761094643e-04, // 220
-1.875475535824517e-02, // 221
-4.982094594654668e+02, // 222
 2.676028686220125e-01, // 223
-9.603967450414284e+02, // 224
 1.814094038045042e+02, // 225
 4.622978572818983e+03, // 226
 1.586888835369008e-04, // 227
-3.238267282004546e-02, // 228
-7.594644056747908e+02, // 229
 3.852313451596073e-09, // 230
-2.497184171637709e+00, // 231
 1.231274709902003e+01, // 232
-4.627756904985868e-04, // 233
-9.317961477556441e-09, // 234
 3.985273846631145e-04, // 235
-3.413176855430123e+02, // 236
 2.974173048739033e+03, // 237
-1.418789826099833e-04, // 238
 1.105583244367092e+01, // 239
 2.336497026713911e+02, // 240
-2.219599876034059e-02, // 241
-1.529689514811186e-03, // 242
 2.971997467261536e+01, // 243
 3.213377986527967e+01, // 244
-1.045622442211491e+01, // 245
 1.243078897941196e+03, // 246
-1.332855703443838e-03, // 247
-4.687681641952115e-02, // 248
-2.233082257137705e+03, // 249
-4.109314504451234e-05, // 250
-2.230180465938499e+01, // 251
 1.726463511673800e-04, // 252
-4.543663445257977e+00, // 253
-6.092354974337531e-02, // 254
 6.748120873157222e-01, // 255
 4.976008111231030e-05, // 256
 8.809954778389600e-01, // 257
 1.020793698797789e+03, // 258
 3.373607645951694e+03, // 259
 7.199455573293006e+02, // 260
 5.081361346376717e+01, // 261
 1.257531367299558e+00, // 262
 6.415456104195287e+03, // 263
 3.987765735535033e+00, // 264
-5.224093721504208e+01, // 265
-6.994826850022373e+02, // 266
-1.497624999457563e+01, // 267
 1.732624762163312e+02, // 268
-2.331295676350790e-04, // 269
-2.044801563877174e-01, // 270
-1.108584158068594e+03, // 271
 2.855773009483748e+03, // 272
-1.800686727009565e-02, // 273
 2.460343632205791e-01, // 274
-1.386529114882643e+03, // 275
-6.379912887686925e-01, // 276
 1.761972919984383e+04, // 277
-4.618703092829962e-09, // 278
 6.387267476354817e+01, // 279
-3.728551632176549e+03, // 280
 2.040879982581382e-02, // 281
 4.487284818922681e+03, // 282
 2.105693164026185e-04, // 283
-3.677040633392725e-03, // 284
-4.400259936804862e+03, // 285
 4.577801472437438e+02, // 286
 6.457420288981935e+00, // 287
-8.388154174327107e-07, // 288
-4.956531275763009e+01, // 289
-8.131521797571200e+00, // 290
-4.093416141263706e+02, // 291
-2.971131283246284e+01, // 292
-2.126865466056073e+01, // 293
-2.157726095081300e+00, // 294
-1.262018658292171e+03, // 295
-3.030205267835228e+02, // 296
-9.537474241681558e-01, // 297
 4.020503116984650e-04, // 298
 1.430343006073042e+01, // 299
-3.424395646159210e+01, // 300
-6.459663521959719e-05, // 301
 9.825917062983344e+03, // 302
-2.160991349562942e-02, // 303
 1.846247673064891e-03, // 304
-1.252603742226546e-11, // 305
 4.710958053299293e-01, // 306
 2.385522385480870e+00, // 307
 3.553186268298606e-02, // 308
-8.057493497265912e+02, // 309
 8.288142297717677e-05, // 310
 3.612855226113974e-01, // 311
-1.143955343285040e+00, // 312
 7.068983172475199e-05, // 313
 5.489784665792775e+00, // 314
 1.107271526861000e-01, // 315
 2.829862436415020e+00, // 316
-2.672932551884699e+03, // 317
 1.436171209876937e+03, // 318
-4.780170250652216e+02, // 319
 9.123160753570115e-06, // 320
-2.342256458101883e-01, // 321
 5.030718741985669e+02, // 322
 2.316357855787135e-03, // 323
 1.961640443347234e+03, // 324
-7.847470296349539e+00, // 325
-1.424398592629256e+00, // 326
-1.019238367729599e-02, // 327
 7.501396785985195e+00, // 328
-3.066954633048206e-06, // 329
-2.213597341132716e+01, // 330
 4.229154143277857e-01, // 331
 5.603053896266793e+03, // 332
-1.206154198074799e-06, // 333
 2.091227673441703e+03, // 334
 5.718493874193080e+03, // 335
 1.693848093187701e+02, // 336
 4.557735398383355e+03, // 337
 6.825236517532907e+01, // 338
 6.857214206151257e-04, // 339
-1.389715763831038e-02, // 340
-2.239145461440803e+03, // 341
 1.277046899982001e-05, // 342
 5.523506793836701e+01, // 343
 3.452034813876273e-04, // 344
-5.852815545346799e-02, // 345
-7.954593673562969e+03, // 346
-1.339287195202207e-05, // 347
 5.263432225522903e+00, // 348
-1.227953221155687e+02, // 349
-1.405426339310303e+00, // 350
 7.787262420826561e-01, // 351
 4.473003125606279e-09, // 352
 1.094325032251344e-04, // 353
 5.916235652845430e+00, // 354
-8.552994848164856e+02, // 355
-2.432727662689261e+03, // 356
 3.673306044599970e-05, // 357
 1.708565016199652e+02, // 358
 2.088404666775530e+03, // 359
 5.423024098534728e-07, // 360
-2.462632895706893e+00, // 361
-7.773465309256761e+03, // 362
 5.759605609683924e+01, // 363
 3.259697401926016e+03, // 364
 4.168437140034587e+03, // 365
-4.360736575662389e+03, // 366
 4.150227036503358e+03, // 367
 3.470671225207984e-04, // 368
-3.763101306565095e+01, // 369
-6.258847618943072e+00, // 370
-7.876916717127198e+02, // 371
-3.641196918470724e+00, // 372
-1.611704127222041e-04, // 373
-4.544361508884036e+03, // 374
-8.362004955323879e-04, // 375
-4.043188121366003e+03, // 376
 7.989398878530898e-05, // 377
 2.083487824002359e+00, // 378
 5.136269371865207e+01, // 379
-3.765221500352277e-06, // 380
 6.134649980821239e+02, // 381
 1.525531219311751e-03, // 382
 1.811909087450972e+01, // 383
-1.665072592094201e-07, // 384
-1.690766154248622e-03, // 385
 5.279968656873849e+01, // 386
-3.346744128257385e-06, // 387
-3.701002521366293e-01, // 388
-2.033952777751174e-05, // 389
 3.425034593671228e+01, // 390
 4.974425844199276e-04, // 391
-2.920318795411848e+00, // 392
 6.994166954902586e-04, // 393
-4.210213725195006e+02, // 394
-9.722070612800866e+01, // 395
 1.234496309539675e+02, // 396
 2.521370747494897e-06, // 397
 1.778318302252585e+02, // 398
-2.954167614360464e-04, // 399
-9.388470883518377e+01, // 400
-4.430937535929163e+03, // 401
 1.751981919631373e-03, // 402
-4.974464119565554e+03, // 403
 7.671792965850829e-02, // 404
-1.161759473166657e+00, // 405
 1.621548926054810e+00, // 406
 4.750344959055921e+02, // 407
-9.212362147360045e+01, // 408
 8.000480967670871e-02, // 409
 3.179137326130189e-03, // 410
-4.172923251281773e-03, // 411
-1.438175858833355e+02, // 412
 2.064770212372089e+00, // 413
 2.455432682219075e-03, // 414
 1.096833001434654e+00, // 415
-7.085612207209273e-02, // 416
-2.699580026975488e+00, // 417
 4.517782171630089e+03, // 418
 7.353314402986603e+00, // 419
-2.295168991476206e-01, // 420
 1.556115324470050e-01, // 421
 5.059761755467955e+03, // 422
-2.561380286022736e-03, // 423
-1.803011518639141e+03, // 424
 5.379203007005531e-09, // 425
-2.115138928608214e+01, // 426
 9.982877301118462e-05, // 427
 1.388492939753526e+01, // 428
-1.941730176645402e+03, // 429
-1.069705325888303e+04, // 430
-1.115966319948977e-06, // 431
-1.641577495563202e+00, // 432
-1.405979725833772e-04, // 433
 9.244898971688168e-06, // 434
-2.244758593785686e+03, // 435
-6.084896770061300e+02, // 436
-6.519431512285841e+03, // 437
-3.892684915659404e+03, // 438
-2.414575338642191e-01, // 439
 9.747968598817413e-01, // 440
-8.792912355278726e+03, // 441
-4.373205623452554e+00, // 442
-1.871824390878744e+00, // 443
 2.158049103636035e-08, // 444
-4.483039727167173e-04, // 445
-1.736870375157641e+00, // 446
 2.143721762243272e-06, // 447
 6.780374401863984e+03, // 448
-1.379659666498807e-06, // 449
-1.228756606170186e-06, // 450
-1.154823629008868e+03, // 451
 9.068296431829507e+02, // 452
-5.998731507759092e-03, // 453
 1.920844546962107e+03, // 454
-2.440364338675749e+01, // 455
 2.972554558018558e+02, // 456
 2.210771097859394e+03, // 457
-2.777904997131138e-05, // 458
 3.495152817617078e+02, // 459
-6.792229684146315e-01, // 460
-1.551570888923184e-04, // 461
 1.934425612217051e-03, // 462
 2.203181670493765e-02, // 463
-1.523622249631565e-02, // 464
-2.267273877064825e+03, // 465
-1.008114268817242e+02, // 466
-1.178842029943556e-01, // 467
 3.971996073489651e-07, // 468
-4.286920503568187e+03, // 469
-5.855956908926249e-02, // 470
 2.696897777246322e+00, // 471
 2.363721239388202e-01, // 472
 7.884652500624035e+03, // 473
 6.058254986227661e+03, // 474
 5.089546702973281e+01, // 475
 7.567863761110945e+03, // 476
-4.413504739712962e+03, // 477
-1.068163836926896e-02, // 478
 3.461317903820922e-04, // 479
 3.228634120150262e+03, // 480
 9.889017955998427e+02, // 481
-1.307734606786301e-01, // 482
 1.038253681584437e+03, // 483
 8.482857886888497e+01, // 484
-1.426716694195997e-03, // 485
-4.278257301060693e+03, // 486
-5.968298229513981e-04, // 487
 2.107942835491121e+03, // 488
 2.374695762477320e-06, // 489
 1.559500031190763e-03, // 490
-2.458791715001335e-01, // 491
 3.419782690895735e+01, // 492
-4.718420364994754e+03, // 493
 3.479321305295454e-02, // 494
-5.465421243206745e+00, // 495
 1.379977602740861e+03, // 496
 1.827612072626021e+03, // 497
 4.853479611830429e-04, // 498
-1.861497967903791e+01, // 499
 3.188116961975228e-05, // 500
 9.688156895029992e+02, // 501
 3.161376403194486e-01, // 502
-1.562229994536345e-03, // 503
 6.950326466920707e-05, // 504
 4.928090208382612e+02, // 505
 1.142491676979067e-02, // 506
 4.553852200082209e+03, // 507
-6.642140125119847e-02, // 508
 7.656081386993519e+03, // 509
-2.364318096025502e+03, // 510
-2.070693875627090e-08, // 511
 1.473202446422395e+01, // 512
-1.309057900639590e+00, // 513
-5.323731092011824e+03, // 514
-1.267574598272690e+01, // 515
-5.505921760586266e+02, // 516
 1.657570169133386e+03, // 517
 7.649745697283516e-06, // 518
 3.109213413078699e-04, // 519
 8.392466434955956e-02, // 520
-5.873557749284644e-02, // 521
 1.231950306204390e-03, // 522
-8.408899694638348e-02, // 523
 8.212085460664011e+03, // 524
 1.961496268616506e-02, // 525
-2.833915164692006e-07, // 526
 1.732597868579498e+01, // 527
-4.423343141692810e+03, // 528
 1.167191827315269e-05, // 529
 1.261445683822447e+00, // 530
-1.783495208204162e-05, // 531
-1.076387063070184e+01, // 532
-4.488047568644487e-01, // 533
 2.077742677748486e+00, // 534
-1.291972994639717e+02, // 535
-4.983836869435809e-11, // 536
-1.272580696495992e+01, // 537
 1.178374353916251e+03, // 538
 6.296591993031207e-02, // 539
-6.136077312430710e+03, // 540
-2.475861932211187e+03, // 541
-8.438545773209366e+03, // 542
-1.036351040363150e+01, // 543
 1.548161885542939e+01, // 544
 4.767423347776423e+03, // 545
-1.922062197905617e-02, // 546
 1.363532946422873e+00, // 547
 4.064399109452028e+03, // 548
-7.088175850341413e+02, // 549
 2.370477584786778e-01, // 550
-4.520585567989708e-05, // 551
-1.551791613656452e+03, // 552
 2.927156264246796e+01, // 553
-2.894282207705841e+02, // 554
-3.238190162671758e-06, // 555
-3.344641596594280e-04, // 556
 3.019944554512241e-03, // 557
-6.738933860507422e-04, // 558
-1.435558529673189e-08, // 559
 1.038472005934949e+02, // 560
 2.756864969218620e-02, // 561
 9.092213651221705e+01, // 562
 3.092047850921324e+00, // 563
 1.487574375050371e+03, // 564
-3.820672455661318e+03, // 565
-1.282260870007384e+02, // 566
 4.216639257253433e-02, // 567
-1.180652939734566e+00, // 568
 3.608172857075826e+00, // 569
-1.129284434397208e+01, // 570
-3.706631717842190e+03, // 571
 1.028391114305999e+02, // 572
 2.982893912785817e+02, // 573
 1.715348014814463e+01, // 574
 1.007075958086568e+00, // 575
 2.515466143548696e-03, // 576
 2.200778086307747e+01, // 577
-5.757937785056102e+03, // 578
 2.516464099338859e+03, // 579
 4.896007052225945e-06, // 580
 4.302021613789660e+00, // 581
-6.235966998292720e+03, // 582
 3.277405849937205e+01, // 583
-1.564738277730774e+03, // 584
-2.378700019969180e+00, // 585
-6.937795211993624e+03, // 586
-3.683701498607461e+00, // 587
 2.156729982241354e+01, // 588
-3.359950248570078e-02, // 589
-6.720922414338114e+03, // 590
-7.163311817005975e+02, // 591
 1.310655018830682e+04, // 592
-3.381703454927924e+03, // 593
 4.319610018163781e+03, // 594
 1.561004216790050e+04, // 595
-3.816513569645753e+02; // 596

}
