netcdf x1b_A1B4_v1x {
  // global attributes 
  :name = "x1b_A1B4_v1x<4>";
  :d_AB =  3.638311877798190e+00; // A^(-1))
  :k_AB =  1.464018301067568e+00; // A^(-1))
  :d_BB =  5.751244385369464e+00; // A^(-1))
  :k_BB =  1.179948162368445e+00; // A^(-1))
  dimensions:
  poly = 82;
  variables:
    double poly(poly);
data:
poly =
-1.412540410682738e+01, // 0
 6.348071674423490e+01, // 1
-2.494104080014214e-01, // 2
 1.287386017393248e+00, // 3
 1.280936023457195e+00, // 4
-2.476039467134847e-01, // 5
-3.018156930230866e+00, // 6
-1.294171922442718e-01, // 7
-6.694601998362794e+00, // 8
 1.505064324110866e-02, // 9
-7.551000138877534e-02, // 10
-3.216979266518568e-03, // 11
 1.498578835725977e-02, // 12
-3.051251925228073e-03, // 13
 7.113073110317622e-03, // 14
-7.622949770708978e-02, // 15
-3.685028049639309e-02, // 16
 1.492713980978938e-02, // 17
 1.448091463248669e-02, // 18
 1.912288899767240e-01, // 19
-1.370173862460179e-03, // 20
-3.023903616285796e-03, // 21
-3.746858231675752e-02, // 22
-7.529807392146101e-02, // 23
 7.364731060748982e-03, // 24
 3.910473750156533e-01, // 25
-4.548715651419601e-04, // 26
-1.426453832261230e-03, // 27
 5.824662752352389e-02, // 28
-5.136480608917194e-06, // 29
-2.315065848485741e-05, // 30
-3.852662729904995e-06, // 31
 4.793286016461522e-05, // 32
 1.040822462593905e-04, // 33
-9.820390188456134e-06, // 34
 5.024145741536724e-05, // 35
 4.999526902547422e-05, // 36
 1.191253241717275e-03, // 37
 3.805187605503457e-04, // 38
-4.960711696395867e-04, // 39
-2.421223638266793e-04, // 40
-2.319913173120385e-04, // 41
-4.919131337643380e-04, // 42
-4.840194607995541e-04, // 43
-2.420115092667065e-04, // 44
-8.224106865365000e-07, // 45
-1.138844047628821e-04, // 46
-9.970969904961424e-06, // 47
 5.060079935499033e-05, // 48
-2.461880351912312e-04, // 49
-2.442403954985514e-04, // 50
-1.017771908283941e-05, // 51
-2.373305653197363e-04, // 52
 4.969581732030054e-05, // 53
 1.746543876588412e-05, // 54
 1.188582429443428e-03, // 55
-2.197198754686991e-05, // 56
-1.012226346030958e-05, // 57
-2.499549722695699e-04, // 58
-1.894234601867977e-03, // 59
 2.419928607107403e-03, // 60
 4.810318219735285e-05, // 61
 1.028030134871160e-04, // 62
 1.202343559257283e-03, // 63
-4.947518311046871e-04, // 64
 1.799753304148982e-05, // 65
-3.800783595536632e-06, // 66
-2.975574781864015e-03, // 67
 1.021702528624513e-04, // 68
 1.207763034616611e-03, // 69
-4.844611416628889e-04, // 70
 1.067922523814582e-04, // 71
-6.053315437023697e-03, // 72
-3.856943832213453e-04, // 73
 3.656909073640143e-04, // 74
 2.452343573050680e-03, // 75
-1.187970518323738e-04, // 76
 1.019309601749661e-04, // 77
-5.007816061989860e-04, // 78
-5.539141268590202e-06, // 79
-1.214349481166761e-02, // 80
 9.586566907261393e-05; // 81

}
