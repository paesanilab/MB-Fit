netcdf x2b_A1B2_A1B2_v1x {
  // global attributes 
  :name = "x2b_A1B2_A1B2_v1x<3>";
  :d_intra_AB =  2.999999994687844e+00; // A^(-1))
  :k_intra_AB =  1.897121755696661e+00; // A^(-1))
  :d_intra_BB =  2.733301180397604e+00; // A^(-1))
  :k_intra_BB =  1.999964905871657e+00; // A^(-1))
  :d_AA =  6.999988545419143e+00; // A^(-1))
  :k_AA =  1.118155783780181e+00; // A^(-1))
  :d_AB =  2.525251147612977e+00; // A^(-1))
  :k_AB =  2.250483599544201e+00; // A^(-1))
  :d_BB =  3.369112299819810e+00; // A^(-1))
  :k_BB =  1.869098220328727e+00; // A^(-1))
  :r2i =  6.000000000000000e+00; // A
  :r2f =  7.000000000000000e+00; // A
  dimensions:
  poly = 134;
  variables:
    double poly(poly);
data:
poly =
 7.692545786871643e-01, // 0
-1.248026521860368e+00, // 1
 1.133017547512339e-01, // 2
 1.062026246780831e+00, // 3
-4.460232101603538e+01, // 4
-5.727165413283573e+01, // 5
 3.945796780580039e+01, // 6
-2.882420552278039e+00, // 7
 2.930396981328015e-01, // 8
 2.691714223861724e+00, // 9
 5.435890073868101e+01, // 10
-6.926013511565102e+01, // 11
-3.286525609024367e+02, // 12
-1.783428573519093e+02, // 13
 8.420721749910154e+00, // 14
-1.730868210137381e+02, // 15
 1.091537252481564e+02, // 16
-1.916412315551173e+01, // 17
 6.097763473248847e-01, // 18
 1.425588661018935e+00, // 19
 1.379566869084238e+01, // 20
-1.843373447360935e+01, // 21
-9.396200114696950e+01, // 22
 4.089103028605907e+01, // 23
-8.772780355116687e-04, // 24
-2.317477942032465e+02, // 25
 3.765855157367505e-04, // 26
-1.451504464786583e+01, // 27
-1.431775504198217e+01, // 28
-2.819111963537485e+02, // 29
 1.790653832971696e+02, // 30
-6.529967498078959e+00, // 31
-3.330259098921666e+01, // 32
-2.670262423400096e+01, // 33
-7.686634371159881e+00, // 34
 9.748307904913506e-06, // 35
-7.996002638691966e+00, // 36
-8.373456934562613e-03, // 37
 2.577590694893530e+01, // 38
 1.641581534051706e+02, // 39
 4.222916443749602e+01, // 40
-6.226064212246886e+00, // 41
 7.038331048109634e+00, // 42
 8.701456439084401e-04, // 43
 8.208036070738819e+02, // 44
 9.046176975837015e+01, // 45
-2.750500771323133e+02, // 46
-5.930297207474858e+00, // 47
 4.295653086262778e+02, // 48
 8.173569646727992e+02, // 49
 7.980028037489499e-04, // 50
-2.318862899601509e+02, // 51
-6.659638463284091e-03, // 52
-6.506218350139274e+01, // 53
 5.667842133279789e-02, // 54
 1.864642766854766e+00, // 55
 6.598807710237890e+01, // 56
 4.410606771621061e+02, // 57
-3.811117734293334e+01, // 58
-9.498028025082722e-06, // 59
 7.407978022854998e-02, // 60
 2.174034367138594e+01, // 61
-4.460960952347717e+01, // 62
 2.166664458381032e+01, // 63
 1.476293155779488e+01, // 64
 6.972194037020004e+00, // 65
-2.080882469137249e-02, // 66
-7.074346027703482e-04, // 67
 2.034828502464065e+02, // 68
-1.398120227018753e+03, // 69
-8.324399685696586e+01, // 70
 5.335863350485933e+00, // 71
-6.577368950204490e+00, // 72
-1.532478589447387e-02, // 73
-3.167963270270458e+02, // 74
-1.647146761238435e+01, // 75
 2.647071350678139e+02, // 76
-7.366965713360072e+00, // 77
 1.323821147276196e-02, // 78
-1.278146703389179e-03, // 79
-4.753649576583515e+00, // 80
-1.254016582644702e+02, // 81
 1.861870517508423e-03, // 82
 4.489780723166075e+02, // 83
-2.872969274200737e-03, // 84
 7.373343156618535e+01, // 85
-7.970736136694589e+01, // 86
 1.067083439491251e-05, // 87
 1.024976839364850e+01, // 88
-7.672961016613841e-06, // 89
 5.285760091871231e+02, // 90
-2.048361416467215e-02, // 91
-7.178829402904340e+01, // 92
 1.076982286410779e+02, // 93
 2.092637327816537e+00, // 94
 2.564061729860584e-01, // 95
 6.962744176902507e+01, // 96
 4.577163190855482e+02, // 97
-1.773219814317316e+02, // 98
 2.260481047456934e-02, // 99
-3.244150191270427e+00, // 100
-1.216185941740856e+02, // 101
 9.840909024697789e+02, // 102
-3.050788750167611e-06, // 103
-1.196218080203027e-03, // 104
-4.323934365206987e+02, // 105
 3.618943703371209e+01, // 106
-3.545765636894432e+01, // 107
 3.654362666428817e-03, // 108
 1.246181187066677e-04, // 109
-4.321596092865234e+01, // 110
 7.945595089574544e+00, // 111
 1.689482250235006e+00, // 112
 4.361858635320031e+02, // 113
-8.249193503434666e-01, // 114
-2.622292157224584e+01, // 115
 9.710823398772929e+00, // 116
 2.292197200564770e+01, // 117
 1.745200534638798e-03, // 118
 1.189644829443358e+02, // 119
-1.576717742038122e+00, // 120
 2.671668941991338e-01, // 121
-1.303757261080900e-03, // 122
-1.585502156992806e-03, // 123
 3.952591414251743e+00, // 124
 2.058404828436811e+00, // 125
 1.710199782583881e-02, // 126
 2.063221348987487e+02, // 127
-7.683290402333907e+01, // 128
-1.291585259477441e+01, // 129
-5.590339658721076e-03, // 130
 7.841024137476606e+01, // 131
 3.333351251960857e-04, // 132
 1.158440768963588e-06; // 133

}
