netcdf x2b_A1B2Z2_D1E2_v1x {
  // global attributes 
  :name = "x2b_A1B2Z2_D1E2_v1x<3>";
  :d_intra_AB =  1.425395556923652e+00; // A^(-1))
  :k_intra_AB =  7.557849235626799e-01; // A^(-1))
  :d_intra_BB =  3.409039281964786e-01; // A^(-1))
  :k_intra_BB =  8.166999895203393e-01; // A^(-1))
  :d_intra_DE =  1.481985906363458e+00; // A^(-1))
  :k_intra_DE =  1.457391527228705e+00; // A^(-1))
  :d_intra_EE =  2.254829240150205e-01; // A^(-1))
  :k_intra_EE =  1.601839361526929e+00; // A^(-1))
  :d_AD =  2.944050311550521e-01; // A^(-1))
  :k_AD =  2.061184634483040e+00; // A^(-1))
  :d_AE =  4.165852882045253e-01; // A^(-1))
  :k_AE =  1.274218490940620e+00; // A^(-1))
  :d_BD =  6.494971448786078e+00; // A^(-1))
  :k_BD =  1.129969995529377e+00; // A^(-1))
  :d_BE =  6.623484503302483e+00; // A^(-1))
  :k_BE =  3.204527815433465e-01; // A^(-1))
  :d_DZ =  2.940735366633505e+00; // A^(-1))
  :k_DZ =  8.566106785352392e-01; // A^(-1))
  :d_EZ =  3.871645863573833e+00; // A^(-1))
  :k_EZ =  1.417544672460083e+00; // A^(-1))
  :r2i =  6.000000000000000e+00; // A
  :r2f =  7.000000000000000e+00; // A
  dimensions:
  poly = 492;
  variables:
    double poly(poly);
data:
poly =
 0.000000000000000e+00, // 0
 0.000000000000000e+00, // 1
 0.000000000000000e+00, // 2
 0.000000000000000e+00, // 3
 0.000000000000000e+00, // 4
 0.000000000000000e+00, // 5
 0.000000000000000e+00, // 6
 0.000000000000000e+00, // 7
 0.000000000000000e+00, // 8
 0.000000000000000e+00, // 9
 0.000000000000000e+00, // 10
 0.000000000000000e+00, // 11
 0.000000000000000e+00, // 12
 0.000000000000000e+00, // 13
 0.000000000000000e+00, // 14
 0.000000000000000e+00, // 15
 0.000000000000000e+00, // 16
 0.000000000000000e+00, // 17
 0.000000000000000e+00, // 18
 0.000000000000000e+00, // 19
 0.000000000000000e+00, // 20
 0.000000000000000e+00, // 21
 0.000000000000000e+00, // 22
 0.000000000000000e+00, // 23
 0.000000000000000e+00, // 24
 0.000000000000000e+00, // 25
 0.000000000000000e+00, // 26
 0.000000000000000e+00, // 27
 0.000000000000000e+00, // 28
 0.000000000000000e+00, // 29
 0.000000000000000e+00, // 30
 0.000000000000000e+00, // 31
 0.000000000000000e+00, // 32
 0.000000000000000e+00, // 33
 0.000000000000000e+00, // 34
 0.000000000000000e+00, // 35
 0.000000000000000e+00, // 36
 0.000000000000000e+00, // 37
 0.000000000000000e+00, // 38
 0.000000000000000e+00, // 39
 0.000000000000000e+00, // 40
 0.000000000000000e+00, // 41
 0.000000000000000e+00, // 42
 0.000000000000000e+00, // 43
 0.000000000000000e+00, // 44
 0.000000000000000e+00, // 45
 0.000000000000000e+00, // 46
 0.000000000000000e+00, // 47
 0.000000000000000e+00, // 48
 0.000000000000000e+00, // 49
 0.000000000000000e+00, // 50
 0.000000000000000e+00, // 51
 0.000000000000000e+00, // 52
 0.000000000000000e+00, // 53
 0.000000000000000e+00, // 54
 0.000000000000000e+00, // 55
 0.000000000000000e+00, // 56
 0.000000000000000e+00, // 57
 0.000000000000000e+00, // 58
 0.000000000000000e+00, // 59
 0.000000000000000e+00, // 60
 0.000000000000000e+00, // 61
 0.000000000000000e+00, // 62
 0.000000000000000e+00, // 63
 0.000000000000000e+00, // 64
 0.000000000000000e+00, // 65
 0.000000000000000e+00, // 66
 0.000000000000000e+00, // 67
 0.000000000000000e+00, // 68
 0.000000000000000e+00, // 69
 0.000000000000000e+00, // 70
 0.000000000000000e+00, // 71
 0.000000000000000e+00, // 72
 0.000000000000000e+00, // 73
 0.000000000000000e+00, // 74
 0.000000000000000e+00, // 75
 0.000000000000000e+00, // 76
 0.000000000000000e+00, // 77
 0.000000000000000e+00, // 78
 0.000000000000000e+00, // 79
 0.000000000000000e+00, // 80
 0.000000000000000e+00, // 81
 0.000000000000000e+00, // 82
 0.000000000000000e+00, // 83
 0.000000000000000e+00, // 84
 0.000000000000000e+00, // 85
 0.000000000000000e+00, // 86
 0.000000000000000e+00, // 87
 0.000000000000000e+00, // 88
 0.000000000000000e+00, // 89
 0.000000000000000e+00, // 90
 0.000000000000000e+00, // 91
 0.000000000000000e+00, // 92
 0.000000000000000e+00, // 93
 0.000000000000000e+00, // 94
 0.000000000000000e+00, // 95
 0.000000000000000e+00, // 96
 0.000000000000000e+00, // 97
 0.000000000000000e+00, // 98
 0.000000000000000e+00, // 99
 0.000000000000000e+00, // 100
 0.000000000000000e+00, // 101
 0.000000000000000e+00, // 102
 0.000000000000000e+00, // 103
 0.000000000000000e+00, // 104
 0.000000000000000e+00, // 105
 0.000000000000000e+00, // 106
 0.000000000000000e+00, // 107
 0.000000000000000e+00, // 108
 0.000000000000000e+00, // 109
 0.000000000000000e+00, // 110
 0.000000000000000e+00, // 111
 0.000000000000000e+00, // 112
 0.000000000000000e+00, // 113
 0.000000000000000e+00, // 114
 0.000000000000000e+00, // 115
 0.000000000000000e+00, // 116
 0.000000000000000e+00, // 117
 0.000000000000000e+00, // 118
 0.000000000000000e+00, // 119
 0.000000000000000e+00, // 120
 0.000000000000000e+00, // 121
 0.000000000000000e+00, // 122
 0.000000000000000e+00, // 123
 0.000000000000000e+00, // 124
 0.000000000000000e+00, // 125
 0.000000000000000e+00, // 126
 0.000000000000000e+00, // 127
 0.000000000000000e+00, // 128
 0.000000000000000e+00, // 129
 0.000000000000000e+00, // 130
 0.000000000000000e+00, // 131
 0.000000000000000e+00, // 132
 0.000000000000000e+00, // 133
 0.000000000000000e+00, // 134
 0.000000000000000e+00, // 135
 0.000000000000000e+00, // 136
 0.000000000000000e+00, // 137
 0.000000000000000e+00, // 138
 0.000000000000000e+00, // 139
 0.000000000000000e+00, // 140
 0.000000000000000e+00, // 141
 0.000000000000000e+00, // 142
 0.000000000000000e+00, // 143
 0.000000000000000e+00, // 144
 0.000000000000000e+00, // 145
 0.000000000000000e+00, // 146
 0.000000000000000e+00, // 147
 0.000000000000000e+00, // 148
 0.000000000000000e+00, // 149
 0.000000000000000e+00, // 150
 0.000000000000000e+00, // 151
 0.000000000000000e+00, // 152
 0.000000000000000e+00, // 153
 0.000000000000000e+00, // 154
 0.000000000000000e+00, // 155
 0.000000000000000e+00, // 156
 0.000000000000000e+00, // 157
 0.000000000000000e+00, // 158
 0.000000000000000e+00, // 159
 0.000000000000000e+00, // 160
 0.000000000000000e+00, // 161
 0.000000000000000e+00, // 162
 0.000000000000000e+00, // 163
 0.000000000000000e+00, // 164
 0.000000000000000e+00, // 165
 0.000000000000000e+00, // 166
 0.000000000000000e+00, // 167
 0.000000000000000e+00, // 168
 0.000000000000000e+00, // 169
 0.000000000000000e+00, // 170
 0.000000000000000e+00, // 171
 0.000000000000000e+00, // 172
 0.000000000000000e+00, // 173
 0.000000000000000e+00, // 174
 0.000000000000000e+00, // 175
 0.000000000000000e+00, // 176
 0.000000000000000e+00, // 177
 0.000000000000000e+00, // 178
 0.000000000000000e+00, // 179
 0.000000000000000e+00, // 180
 0.000000000000000e+00, // 181
 0.000000000000000e+00, // 182
 0.000000000000000e+00, // 183
 0.000000000000000e+00, // 184
 0.000000000000000e+00, // 185
 0.000000000000000e+00, // 186
 0.000000000000000e+00, // 187
 0.000000000000000e+00, // 188
 0.000000000000000e+00, // 189
 0.000000000000000e+00, // 190
 0.000000000000000e+00, // 191
 0.000000000000000e+00, // 192
 0.000000000000000e+00, // 193
 0.000000000000000e+00, // 194
 0.000000000000000e+00, // 195
 0.000000000000000e+00, // 196
 0.000000000000000e+00, // 197
 0.000000000000000e+00, // 198
 0.000000000000000e+00, // 199
 0.000000000000000e+00, // 200
 0.000000000000000e+00, // 201
 0.000000000000000e+00, // 202
 0.000000000000000e+00, // 203
 0.000000000000000e+00, // 204
 0.000000000000000e+00, // 205
 0.000000000000000e+00, // 206
 0.000000000000000e+00, // 207
 0.000000000000000e+00, // 208
 0.000000000000000e+00, // 209
 0.000000000000000e+00, // 210
 0.000000000000000e+00, // 211
 0.000000000000000e+00, // 212
 0.000000000000000e+00, // 213
 0.000000000000000e+00, // 214
 0.000000000000000e+00, // 215
 0.000000000000000e+00, // 216
 0.000000000000000e+00, // 217
 0.000000000000000e+00, // 218
 0.000000000000000e+00, // 219
 0.000000000000000e+00, // 220
 0.000000000000000e+00, // 221
 0.000000000000000e+00, // 222
 0.000000000000000e+00, // 223
 0.000000000000000e+00, // 224
 0.000000000000000e+00, // 225
 0.000000000000000e+00, // 226
 0.000000000000000e+00, // 227
 0.000000000000000e+00, // 228
 0.000000000000000e+00, // 229
 0.000000000000000e+00, // 230
 0.000000000000000e+00, // 231
 0.000000000000000e+00, // 232
 0.000000000000000e+00, // 233
 0.000000000000000e+00, // 234
 0.000000000000000e+00, // 235
 0.000000000000000e+00, // 236
 0.000000000000000e+00, // 237
 0.000000000000000e+00, // 238
 0.000000000000000e+00, // 239
 0.000000000000000e+00, // 240
 0.000000000000000e+00, // 241
 0.000000000000000e+00, // 242
 0.000000000000000e+00, // 243
 0.000000000000000e+00, // 244
 0.000000000000000e+00, // 245
 0.000000000000000e+00, // 246
 0.000000000000000e+00, // 247
 0.000000000000000e+00, // 248
 0.000000000000000e+00, // 249
 0.000000000000000e+00, // 250
 0.000000000000000e+00, // 251
 0.000000000000000e+00, // 252
 0.000000000000000e+00, // 253
 0.000000000000000e+00, // 254
 0.000000000000000e+00, // 255
 0.000000000000000e+00, // 256
 0.000000000000000e+00, // 257
 0.000000000000000e+00, // 258
 0.000000000000000e+00, // 259
 0.000000000000000e+00, // 260
 0.000000000000000e+00, // 261
 0.000000000000000e+00, // 262
 0.000000000000000e+00, // 263
 0.000000000000000e+00, // 264
 0.000000000000000e+00, // 265
 0.000000000000000e+00, // 266
 0.000000000000000e+00, // 267
 0.000000000000000e+00, // 268
 0.000000000000000e+00, // 269
 0.000000000000000e+00, // 270
 0.000000000000000e+00, // 271
 0.000000000000000e+00, // 272
 0.000000000000000e+00, // 273
 0.000000000000000e+00, // 274
 0.000000000000000e+00, // 275
 0.000000000000000e+00, // 276
 0.000000000000000e+00, // 277
 0.000000000000000e+00, // 278
 0.000000000000000e+00, // 279
 0.000000000000000e+00, // 280
 0.000000000000000e+00, // 281
 0.000000000000000e+00, // 282
 0.000000000000000e+00, // 283
 0.000000000000000e+00, // 284
 0.000000000000000e+00, // 285
 0.000000000000000e+00, // 286
 0.000000000000000e+00, // 287
 0.000000000000000e+00, // 288
 0.000000000000000e+00, // 289
 0.000000000000000e+00, // 290
 0.000000000000000e+00, // 291
 0.000000000000000e+00, // 292
 0.000000000000000e+00, // 293
 0.000000000000000e+00, // 294
 0.000000000000000e+00, // 295
 0.000000000000000e+00, // 296
 0.000000000000000e+00, // 297
 0.000000000000000e+00, // 298
 0.000000000000000e+00, // 299
 0.000000000000000e+00, // 300
 0.000000000000000e+00, // 301
 0.000000000000000e+00, // 302
 0.000000000000000e+00, // 303
 0.000000000000000e+00, // 304
 0.000000000000000e+00, // 305
 0.000000000000000e+00, // 306
 0.000000000000000e+00, // 307
 0.000000000000000e+00, // 308
 0.000000000000000e+00, // 309
 0.000000000000000e+00, // 310
 0.000000000000000e+00, // 311
 0.000000000000000e+00, // 312
 0.000000000000000e+00, // 313
 0.000000000000000e+00, // 314
 0.000000000000000e+00, // 315
 0.000000000000000e+00, // 316
 0.000000000000000e+00, // 317
 0.000000000000000e+00, // 318
 0.000000000000000e+00, // 319
 0.000000000000000e+00, // 320
 0.000000000000000e+00, // 321
 0.000000000000000e+00, // 322
 0.000000000000000e+00, // 323
 0.000000000000000e+00, // 324
 0.000000000000000e+00, // 325
 0.000000000000000e+00, // 326
 0.000000000000000e+00, // 327
 0.000000000000000e+00, // 328
 0.000000000000000e+00, // 329
 0.000000000000000e+00, // 330
 0.000000000000000e+00, // 331
 0.000000000000000e+00, // 332
 0.000000000000000e+00, // 333
 0.000000000000000e+00, // 334
 0.000000000000000e+00, // 335
 0.000000000000000e+00, // 336
 0.000000000000000e+00, // 337
 0.000000000000000e+00, // 338
 0.000000000000000e+00, // 339
 0.000000000000000e+00, // 340
 0.000000000000000e+00, // 341
 0.000000000000000e+00, // 342
 0.000000000000000e+00, // 343
 0.000000000000000e+00, // 344
 0.000000000000000e+00, // 345
 0.000000000000000e+00, // 346
 0.000000000000000e+00, // 347
 0.000000000000000e+00, // 348
 0.000000000000000e+00, // 349
 0.000000000000000e+00, // 350
 0.000000000000000e+00, // 351
 0.000000000000000e+00, // 352
 0.000000000000000e+00, // 353
 0.000000000000000e+00, // 354
 0.000000000000000e+00, // 355
 0.000000000000000e+00, // 356
 0.000000000000000e+00, // 357
 0.000000000000000e+00, // 358
 0.000000000000000e+00, // 359
 0.000000000000000e+00, // 360
 0.000000000000000e+00, // 361
 0.000000000000000e+00, // 362
 0.000000000000000e+00, // 363
 0.000000000000000e+00, // 364
 0.000000000000000e+00, // 365
 0.000000000000000e+00, // 366
 0.000000000000000e+00, // 367
 0.000000000000000e+00, // 368
 0.000000000000000e+00, // 369
 0.000000000000000e+00, // 370
 0.000000000000000e+00, // 371
 0.000000000000000e+00, // 372
 0.000000000000000e+00, // 373
 0.000000000000000e+00, // 374
 0.000000000000000e+00, // 375
 0.000000000000000e+00, // 376
 0.000000000000000e+00, // 377
 0.000000000000000e+00, // 378
 0.000000000000000e+00, // 379
 0.000000000000000e+00, // 380
 0.000000000000000e+00, // 381
 0.000000000000000e+00, // 382
 0.000000000000000e+00, // 383
 0.000000000000000e+00, // 384
 0.000000000000000e+00, // 385
 0.000000000000000e+00, // 386
 0.000000000000000e+00, // 387
 0.000000000000000e+00, // 388
 0.000000000000000e+00, // 389
 0.000000000000000e+00, // 390
 0.000000000000000e+00, // 391
 0.000000000000000e+00, // 392
 0.000000000000000e+00, // 393
 0.000000000000000e+00, // 394
 0.000000000000000e+00, // 395
 0.000000000000000e+00, // 396
 0.000000000000000e+00, // 397
 0.000000000000000e+00, // 398
 0.000000000000000e+00, // 399
 0.000000000000000e+00, // 400
 0.000000000000000e+00, // 401
 0.000000000000000e+00, // 402
 0.000000000000000e+00, // 403
 0.000000000000000e+00, // 404
 0.000000000000000e+00, // 405
 0.000000000000000e+00, // 406
 0.000000000000000e+00, // 407
 0.000000000000000e+00, // 408
 0.000000000000000e+00, // 409
 0.000000000000000e+00, // 410
 0.000000000000000e+00, // 411
 0.000000000000000e+00, // 412
 0.000000000000000e+00, // 413
 0.000000000000000e+00, // 414
 0.000000000000000e+00, // 415
 0.000000000000000e+00, // 416
 0.000000000000000e+00, // 417
 0.000000000000000e+00, // 418
 0.000000000000000e+00, // 419
 0.000000000000000e+00, // 420
 0.000000000000000e+00, // 421
 0.000000000000000e+00, // 422
 0.000000000000000e+00, // 423
 0.000000000000000e+00, // 424
 0.000000000000000e+00, // 425
 0.000000000000000e+00, // 426
 0.000000000000000e+00, // 427
 0.000000000000000e+00, // 428
 0.000000000000000e+00, // 429
 0.000000000000000e+00, // 430
 0.000000000000000e+00, // 431
 0.000000000000000e+00, // 432
 0.000000000000000e+00, // 433
 0.000000000000000e+00, // 434
 0.000000000000000e+00, // 435
 0.000000000000000e+00, // 436
 0.000000000000000e+00, // 437
 0.000000000000000e+00, // 438
 0.000000000000000e+00, // 439
 0.000000000000000e+00, // 440
 0.000000000000000e+00, // 441
 0.000000000000000e+00, // 442
 0.000000000000000e+00, // 443
 0.000000000000000e+00, // 444
 0.000000000000000e+00, // 445
 0.000000000000000e+00, // 446
 0.000000000000000e+00, // 447
 0.000000000000000e+00, // 448
 0.000000000000000e+00, // 449
 0.000000000000000e+00, // 450
 0.000000000000000e+00, // 451
 0.000000000000000e+00, // 452
 0.000000000000000e+00, // 453
 0.000000000000000e+00, // 454
 0.000000000000000e+00, // 455
 0.000000000000000e+00, // 456
 0.000000000000000e+00, // 457
 0.000000000000000e+00, // 458
 0.000000000000000e+00, // 459
 0.000000000000000e+00, // 460
 0.000000000000000e+00, // 461
 0.000000000000000e+00, // 462
 0.000000000000000e+00, // 463
 0.000000000000000e+00, // 464
 0.000000000000000e+00, // 465
 0.000000000000000e+00, // 466
 0.000000000000000e+00, // 467
 0.000000000000000e+00, // 468
 0.000000000000000e+00, // 469
 0.000000000000000e+00, // 470
 0.000000000000000e+00, // 471
 0.000000000000000e+00, // 472
 0.000000000000000e+00, // 473
 0.000000000000000e+00, // 474
 0.000000000000000e+00, // 475
 0.000000000000000e+00, // 476
 0.000000000000000e+00, // 477
 0.000000000000000e+00, // 478
 0.000000000000000e+00, // 479
 0.000000000000000e+00, // 480
 0.000000000000000e+00, // 481
 0.000000000000000e+00, // 482
 0.000000000000000e+00, // 483
 0.000000000000000e+00, // 484
 0.000000000000000e+00, // 485
 0.000000000000000e+00, // 486
 0.000000000000000e+00, // 487
 0.000000000000000e+00, // 488
 0.000000000000000e+00, // 489
 0.000000000000000e+00, // 490
 0.000000000000000e+00; // 491

}
