netcdf x2b_A1B2_A1B2_v1x {
  // global attributes 
  :name = "x2b_A1B2_A1B2_v1x<4>";
  :d_intra_AB =  2.999999009415175e+00; // A^(-1))
  :k_intra_AB =  1.927742824782188e+00; // A^(-1))
  :d_intra_BB =  2.847826708059092e+00; // A^(-1))
  :k_intra_BB =  2.842787560401611e-01; // A^(-1))
  :d_AA =  3.968587662548076e+00; // A^(-1))
  :k_AA =  1.219517528031537e+00; // A^(-1))
  :d_AB =  3.279627749122528e+00; // A^(-1))
  :k_AB =  2.033497636561858e+00; // A^(-1))
  :d_BB =  5.001923151566628e+00; // A^(-1))
  :k_BB =  1.237413265348416e+00; // A^(-1))
  :r2i =  6.000000000000000e+00; // A
  :r2f =  7.000000000000000e+00; // A
  dimensions:
  poly = 597;
  variables:
    double poly(poly);
data:
poly =
-1.031207655862965e-03, // 0
 4.995080204928852e-03, // 1
-5.806886972756709e-03, // 2
 3.430096576072369e-03, // 3
 2.630376394101821e+00, // 4
-4.958417055555740e-02, // 5
 4.251967654846953e-01, // 6
 1.326716309614572e-03, // 7
 5.472425461503635e-03, // 8
-7.312980835907776e-02, // 9
-1.310796322261112e-02, // 10
 1.015285238706463e+00, // 11
-4.792450666385015e-01, // 12
 1.303084745196926e-01, // 13
 1.112375731612144e-02, // 14
 2.552710470553624e-01, // 15
-2.816847617454780e-01, // 16
-5.653337622999041e-02, // 17
-4.133687576457991e-03, // 18
 8.300360530800520e-02, // 19
-5.421033338770292e-01, // 20
-6.074637594784896e-02, // 21
 1.317572571967517e-02, // 22
-2.281900823556336e+00, // 23
-9.172078133302294e+01, // 24
 1.567638701977329e+01, // 25
 1.114251388664594e+01, // 26
-8.642110294722397e-01, // 27
 8.661127876027688e-01, // 28
-3.056478437807362e-01, // 29
 1.002566563225861e+00, // 30
 4.505466497370750e+01, // 31
 1.134444570681847e+00, // 32
 3.282633914020949e-01, // 33
 1.432416012446832e-01, // 34
 1.618460718392840e+01, // 35
 8.816602542623984e+00, // 36
-6.821791638231281e+00, // 37
-6.762309200799837e+00, // 38
 9.876057165306451e-01, // 39
-4.955677568174268e-01, // 40
-6.353256229995893e-03, // 41
-2.277819448183229e+00, // 42
-5.860159347651502e+00, // 43
-4.457684551246173e-01, // 44
 2.584374442030949e+00, // 45
-2.753681720916091e-01, // 46
-1.323787264372508e+00, // 47
 2.433683605101399e-01, // 48
-4.279809347058413e-01, // 49
-3.186386398826795e+00, // 50
-2.709958574620638e-01, // 51
 1.075536209897441e+01, // 52
-7.294770575595625e+00, // 53
 2.934392479662556e+01, // 54
 1.547553499019147e-02, // 55
 3.518060845274660e+01, // 56
 2.650645881611058e-01, // 57
 3.146407022548532e+00, // 58
 1.703319791603978e+00, // 59
 3.272307512656807e-03, // 60
-8.607607074086038e+00, // 61
 4.549310605277341e-01, // 62
-2.714809383632388e+00, // 63
-4.512324820814330e+00, // 64
 5.336899899016237e+00, // 65
-1.035762319852744e+01, // 66
-5.116497089033112e+01, // 67
-1.457284735086362e+00, // 68
-1.674652970511178e-01, // 69
-8.341908485549524e+00, // 70
-5.019170597936591e-01, // 71
 4.593202453829964e+01, // 72
-2.351012924193112e+01, // 73
-9.321159682936568e-01, // 74
-1.078431500020082e-01, // 75
-8.785318555978838e+00, // 76
-6.208126879135273e+00, // 77
 5.717219984914811e+01, // 78
-9.673367891365453e-02, // 79
-4.822177941083996e+00, // 80
 7.911422418928747e+00, // 81
 7.956541162013587e+00, // 82
 1.264517034996192e-01, // 83
-9.792291662036474e+00, // 84
-5.621196701491325e-02, // 85
 4.589173636557567e-01, // 86
-4.596001104672187e+01, // 87
 8.977375500912730e+01, // 88
 3.316921569632697e+01, // 89
-9.938980307062877e-01, // 90
-1.364200346307584e+01, // 91
-3.792647406695299e-02, // 92
-3.836483996935634e-02, // 93
-2.217224746172846e+00, // 94
 4.556695841240943e+00, // 95
-8.783634406561632e-01, // 96
 1.356981839777926e-01, // 97
 2.586551615052989e+00, // 98
 2.242127609944094e+00, // 99
-4.868665892396750e-03, // 100
-5.208969981541772e-05, // 101
-1.879127949480219e-01, // 102
-2.043653691676173e+01, // 103
-1.678861702201733e+01, // 104
-1.765493397471752e+01, // 105
 2.384428783213813e-02, // 106
-3.179398474678084e-02, // 107
 3.098118154505929e+00, // 108
 3.387393081312878e+01, // 109
-3.614207638974676e-02, // 110
 4.996000957748518e-01, // 111
-6.503307361590400e-04, // 112
 3.718330992199276e-02, // 113
-1.578342807626573e+02, // 114
 3.247631257297610e+00, // 115
-9.425610084928319e-03, // 116
-6.469797371895987e+00, // 117
 5.903406634155888e+00, // 118
-1.560949378461730e+00, // 119
-2.348500003660993e-03, // 120
-1.770664999705271e-03, // 121
 6.416118864990449e+01, // 122
 2.283430940983602e+01, // 123
 2.148632856888326e-02, // 124
 7.687605864027198e-01, // 125
-1.783409572651716e+01, // 126
-1.092967833601752e+00, // 127
 3.431198383597712e+01, // 128
 5.141627654507444e+00, // 129
 3.921343890186205e+01, // 130
-5.705772185473922e-02, // 131
-4.023287731934596e+01, // 132
-9.376573033640874e+00, // 133
 4.946930497344213e-02, // 134
 6.699917099920999e-02, // 135
-2.540172465940627e-04, // 136
 6.888244867649912e+00, // 137
-1.953170781475734e+00, // 138
 3.042018581768499e-01, // 139
 1.890877407268660e-04, // 140
 5.102833979724038e+01, // 141
 4.883585666825350e-01, // 142
-5.503927547548997e+01, // 143
-5.666586148343030e+01, // 144
-1.119068531668491e+00, // 145
-1.519440078728925e-03, // 146
-1.957941568898906e-04, // 147
-4.778236094152091e+00, // 148
 1.495227321362671e-02, // 149
-4.703773526588924e+00, // 150
-1.883416515495141e+00, // 151
 3.919319528864734e-01, // 152
 4.439517942084401e-01, // 153
-1.830899424207754e-01, // 154
-4.060907030277244e+00, // 155
-4.168485852987223e-01, // 156
 1.634799699381614e+00, // 157
-9.721653638457279e+01, // 158
-2.025688039906248e-02, // 159
-1.445196354209205e-01, // 160
 2.948520918863616e+00, // 161
-2.189416219815526e+00, // 162
-1.633039780244224e-03, // 163
-6.173161305110283e+00, // 164
 1.484925632478420e+02, // 165
 2.997084577753030e-02, // 166
 1.467468419503005e+00, // 167
 4.815028299479657e-01, // 168
-1.349398670971037e-04, // 169
 1.413281761588485e+01, // 170
-1.990880914077569e+00, // 171
 1.229493157803220e-01, // 172
 1.961643561375786e+01, // 173
 9.057358550281557e-01, // 174
-5.457647752598212e-02, // 175
-2.134554155120337e-01, // 176
-1.419699284655039e-03, // 177
-4.865072841538401e+00, // 178
 1.118051332410302e+01, // 179
-1.908368156106577e+01, // 180
-2.399005835628223e+00, // 181
-1.116233902504419e+02, // 182
-6.154888474651971e+00, // 183
 2.459323929732650e-03, // 184
-9.034511455291637e+00, // 185
 7.966020004472913e-01, // 186
-2.686798418760613e-05, // 187
-2.783166004290521e-01, // 188
 8.780395707753946e-01, // 189
 1.541073633385116e+01, // 190
 4.705279939266841e+01, // 191
 1.378596691511110e+00, // 192
-3.161471457831639e-01, // 193
-1.940629206051745e-01, // 194
 2.253402303853951e+01, // 195
-4.249702798123711e-01, // 196
 9.579378392428079e-05, // 197
-5.229445775021095e-01, // 198
 9.788389949864248e+00, // 199
 4.845209662457080e-02, // 200
-3.561472172222055e-05, // 201
-3.737694842016555e+01, // 202
-1.836228145409826e+00, // 203
-1.864572214270521e+00, // 204
 1.080774180387122e+01, // 205
-9.616654219944746e+00, // 206
-2.367199145295279e-05, // 207
 1.428533563722217e+01, // 208
-1.335756301688084e+00, // 209
 1.100614815431716e-01, // 210
 2.049705656992061e-04, // 211
 1.073984223202955e-01, // 212
 4.972138015725696e-01, // 213
 8.589751248642151e-01, // 214
 3.625926059801118e-03, // 215
 1.127214111316197e+00, // 216
-6.293366850601581e+00, // 217
-3.262686846594030e+01, // 218
 5.637260363096443e-02, // 219
 4.993521399899870e-01, // 220
 8.384083654336686e-01, // 221
-4.293612575111640e-01, // 222
-5.898496412543022e-01, // 223
-8.535278339591950e-04, // 224
 5.452342714410009e+00, // 225
 1.123056583234507e+01, // 226
-1.719308789117955e-01, // 227
-1.504666727602648e+01, // 228
 4.149302604487418e+01, // 229
-7.801577284364136e-06, // 230
-1.522103983080871e+01, // 231
 1.259483970523682e+00, // 232
 3.702692552500930e-01, // 233
-9.266237672323778e-06, // 234
 9.020861583380059e+00, // 235
 2.557584455532482e+00, // 236
-4.360332146735770e-01, // 237
 9.921148651076921e-05, // 238
 4.887170171307293e+00, // 239
-1.491991696398527e+02, // 240
-1.976359591257076e+01, // 241
 4.467436553121764e-01, // 242
 5.525468110149288e+01, // 243
-9.270584227056777e-01, // 244
-3.369783433016636e+00, // 245
-1.140234111511870e+01, // 246
 3.233710057907739e-01, // 247
 1.432807603142820e+00, // 248
 2.554897718049471e+00, // 249
 6.943751516153411e-05, // 250
-1.366768087240445e-03, // 251
-3.833331255924174e-01, // 252
 2.433676942194881e-01, // 253
 3.898715095932644e-04, // 254
-1.056207655977718e+00, // 255
-3.820729800981224e-05, // 256
-5.781513174047467e-02, // 257
 4.814370808454816e-03, // 258
 7.302211015161897e+01, // 259
 3.714254423034168e+01, // 260
-1.906995794236074e+01, // 261
-1.462344566172534e-01, // 262
-1.340351925116305e+01, // 263
 3.068877973235403e+00, // 264
-5.107277159534062e+00, // 265
-4.431819770371870e-01, // 266
-5.847140511941800e+00, // 267
 3.693160831283026e+01, // 268
-3.207120417493086e-04, // 269
 7.824220118106287e+00, // 270
 3.361021432424140e-03, // 271
-1.331294989110213e+01, // 272
 5.849601815394776e+00, // 273
-8.882383738284551e-04, // 274
-1.734932200244475e-01, // 275
 1.293738611262111e+00, // 276
-2.415002124236444e+01, // 277
-9.475511948846356e-06, // 278
-5.542664768002848e+00, // 279
 5.117415646154889e-01, // 280
-2.041591541624142e+01, // 281
-5.810736164367728e+00, // 282
-1.734184248241146e-05, // 283
-2.231907956552969e+01, // 284
 1.408615156577647e+01, // 285
-2.168957843370290e+00, // 286
 4.491150547021169e+00, // 287
-1.656629177019283e-04, // 288
 1.077120698907685e+02, // 289
-4.376346937469585e+00, // 290
-1.665651660365189e+01, // 291
-4.070710587259861e-01, // 292
 2.983294480624197e+00, // 293
 1.022351897681059e+01, // 294
 2.462305073853068e+00, // 295
 3.774369781162146e+00, // 296
-3.267918490758631e+01, // 297
-8.945390194288059e-04, // 298
 1.170934440540300e+02, // 299
-5.041192351136658e+00, // 300
-8.270026847320345e+00, // 301
-8.624640509034156e-01, // 302
 2.286115508971341e-06, // 303
 4.963347534171958e-04, // 304
 2.075211169275580e-06, // 305
-3.228167043168820e+01, // 306
 2.838821504970046e+01, // 307
 2.721576886067597e-01, // 308
-5.183637322867342e-02, // 309
-2.304543019254548e-05, // 310
-9.689142109475711e+00, // 311
 1.254146459927151e-01, // 312
-2.516223220963576e-05, // 313
 3.158715288837923e+01, // 314
 1.811895080957274e-04, // 315
 4.784901218400944e+01, // 316
 2.804808431560438e+01, // 317
 1.649643236616921e+00, // 318
 1.044355374860058e+01, // 319
-9.922104252875045e-03, // 320
-2.529653002959220e+00, // 321
-4.608038140957375e+00, // 322
 2.167508609809773e-01, // 323
 5.536549733790474e+00, // 324
-1.565396782359744e+01, // 325
-8.142922557375975e+00, // 326
 3.248579292309410e+01, // 327
 1.127570989370199e+02, // 328
 2.156803669472487e-04, // 329
-7.514506155327628e+01, // 330
 4.674423895429985e+01, // 331
 3.279312000114389e-01, // 332
-7.223703423977382e-05, // 333
 4.454168969023031e+00, // 334
 1.266257023091750e+01, // 335
 3.753649836520763e+01, // 336
 1.583974016100707e+00, // 337
 9.713791168694947e+01, // 338
-2.098635446077777e+00, // 339
 2.709724327776579e-03, // 340
-1.823313494982351e-02, // 341
 2.529375837691330e-04, // 342
-1.379571375545230e+00, // 343
 3.307694079281830e-05, // 344
 5.981870531588071e+01, // 345
 3.477600882039858e+01, // 346
-1.455665951230649e+01, // 347
 4.345132538817291e+00, // 348
 2.902297227504874e+01, // 349
-1.641528977196294e+01, // 350
 2.753534668594031e+01, // 351
-8.835810957817599e-06, // 352
 7.318771281832245e+00, // 353
 7.065974444579341e+00, // 354
-4.723656478675428e-01, // 355
-2.518755704764665e-01, // 356
 2.660124554417079e-01, // 357
-2.385903400327394e+01, // 358
 3.763092451532792e-03, // 359
 3.142446659904541e-05, // 360
 2.991637026219276e+00, // 361
-1.698296014028233e-03, // 362
-2.469935031205115e-01, // 363
 4.834587987300753e-01, // 364
 4.030032863978585e-01, // 365
-1.327683280217554e+01, // 366
-3.328758953075864e+01, // 367
 2.360811029925665e-01, // 368
-5.959799882069587e+00, // 369
 1.227667345901177e-01, // 370
-7.917322495802448e+01, // 371
-9.106840438063880e-01, // 372
-8.062838373413310e-06, // 373
-1.905822692729364e+00, // 374
-8.246910396593561e+00, // 375
-1.456997060847798e+01, // 376
-7.227322038010151e-03, // 377
-7.362040018602380e+00, // 378
 2.193683767217629e+00, // 379
 9.954594544396152e-02, // 380
 3.631253060315975e+01, // 381
 3.918776575851779e-04, // 382
-1.067032461581510e+01, // 383
 1.849840486527010e-05, // 384
 2.475192036941537e-01, // 385
-5.292032037054039e+00, // 386
 9.924822438667034e-02, // 387
 1.535795057262605e+00, // 388
 1.356881655426653e+00, // 389
-1.501859407067921e+02, // 390
-1.389308117476780e-05, // 391
 8.002044860487148e+00, // 392
-1.197872566682568e-03, // 393
 7.925208976047959e+01, // 394
-5.675617348830828e+01, // 395
-1.474525503444885e+00, // 396
-1.576072482908959e+01, // 397
 8.818131217418075e+01, // 398
-1.725349037251687e-01, // 399
-8.257498368729010e+01, // 400
 5.444273330835838e+01, // 401
 2.387149809068184e-04, // 402
-4.346909954025148e+00, // 403
-9.297026597580494e-01, // 404
 2.301271869774597e-01, // 405
-3.405322222709909e-01, // 406
-1.474315799031810e+00, // 407
 3.517222165154660e+00, // 408
-3.661580021262063e-01, // 409
 3.237045278251958e+01, // 410
-1.468106205003896e-01, // 411
-1.606122022644306e+01, // 412
-4.160522136745699e+00, // 413
 7.536736011195980e-05, // 414
 2.593234246851732e-01, // 415
-2.351403145652488e+00, // 416
-4.196807513413370e+01, // 417
 1.857853605735486e-02, // 418
-6.161437170939627e+01, // 419
-3.867927881046320e-01, // 420
 5.263045145815909e+01, // 421
-1.295137491121063e+02, // 422
-3.506124737807024e+00, // 423
 3.714904312444797e+01, // 424
-2.578669906375152e-06, // 425
-6.651163444895158e+00, // 426
-1.338801679493059e-06, // 427
-1.302521891165020e+02, // 428
 1.464351833349739e-02, // 429
-2.002603976083598e-02, // 430
 4.617115210259928e-05, // 431
 4.584769776312021e+00, // 432
-3.779817240771525e-05, // 433
-6.204701816699276e-02, // 434
 1.067400605861134e+00, // 435
-2.631984192317315e+01, // 436
-6.124458079257684e+00, // 437
 8.000831099795195e-01, // 438
 9.195422630222794e+00, // 439
-1.127955027729906e-01, // 440
-7.434392948673852e+01, // 441
 1.273104522560691e-01, // 442
 9.193065908458134e-02, // 443
 1.539862987097335e-05, // 444
-5.776804059876093e-04, // 445
 2.255450116352496e+01, // 446
-1.754536522658706e-05, // 447
 2.981729097584134e+00, // 448
-3.700550934707666e-05, // 449
-1.616342538285024e-05, // 450
-3.380961949044291e-02, // 451
-2.027977006726555e-01, // 452
 1.284724081840699e-04, // 453
 7.205263459990174e+01, // 454
-7.324608346481328e+01, // 455
 4.251001746652106e+00, // 456
 1.798552259699106e+01, // 457
 1.044632938015666e-04, // 458
 1.067458778865314e+01, // 459
-4.236554821835410e+00, // 460
-1.719024630179598e-04, // 461
 1.351403953986449e-01, // 462
-1.415086999786587e+00, // 463
 3.164939315396096e-01, // 464
-1.830156804188072e+01, // 465
 2.904492254469466e+01, // 466
-1.005026467986533e-03, // 467
-8.878688726270401e-07, // 468
-1.530187836007182e+01, // 469
-8.032897582990952e-05, // 470
 4.191932741889305e+00, // 471
-4.569243011157390e-01, // 472
 2.717281749181074e+01, // 473
 6.404071956435162e-03, // 474
 6.768650848544830e+01, // 475
-5.565366276343495e-04, // 476
-2.590911993455757e+00, // 477
 2.889440087286910e-05, // 478
 1.003645990394722e-01, // 479
 3.508140737466487e-01, // 480
-4.326950604635093e-02, // 481
 3.183666862150145e-02, // 482
-8.172748546851692e+01, // 483
-8.230429479336247e+01, // 484
 6.525063116061950e-05, // 485
 2.300536797934703e-02, // 486
-2.379546662274918e-01, // 487
 9.564614935477744e-01, // 488
-1.088650292333963e-05, // 489
 9.224805135532739e-03, // 490
-2.365914209577594e+00, // 491
 6.338593676537867e+01, // 492
 3.364802013945002e+00, // 493
 6.007749308807732e-01, // 494
 5.006083190244792e-01, // 495
 2.487509176141508e+00, // 496
 4.126633700750012e+01, // 497
 9.417987716452992e-01, // 498
-1.563980289604820e+01, // 499
 5.049646681758410e-01, // 500
-1.010866139523336e+00, // 501
 1.327935288331334e+01, // 502
 3.157684151862030e-04, // 503
 7.285483266008547e-05, // 504
 1.401159625463951e-01, // 505
 1.396626112311455e-03, // 506
-3.048410148138356e-02, // 507
 1.359866026535208e+01, // 508
 3.248093733615898e-01, // 509
-9.605295147810355e-01, // 510
-1.311325605996701e-05, // 511
-2.839267079683627e-01, // 512
 6.449766101517614e-01, // 513
 1.736654188631296e-02, // 514
 5.393578458296363e+01, // 515
 6.275474762321757e+01, // 516
 1.210943338435102e-01, // 517
-8.413295045531122e-06, // 518
-1.228607462158939e-04, // 519
 1.184331910804888e+01, // 520
-1.270347269331055e+01, // 521
-9.617818170145854e-05, // 522
 1.509369267764597e+01, // 523
 3.134504742014008e-02, // 524
-1.534377875599687e+00, // 525
 8.034445724929603e-06, // 526
 2.581374417768561e+01, // 527
-2.381696670798019e+01, // 528
 4.431493665319849e-01, // 529
 4.717538354290226e-01, // 530
-1.616610539481838e-04, // 531
-5.131211611810218e+00, // 532
-1.097458429083981e+00, // 533
 2.504210721139537e+00, // 534
-1.295185776564562e+02, // 535
 1.717051011165495e-06, // 536
 5.445456768119541e+01, // 537
-7.363332058228332e-02, // 538
 1.419872642984520e-01, // 539
-4.578987392298783e-02, // 540
-3.981428338075813e+01, // 541
 6.501554686091094e-03, // 542
 2.452611500519664e+00, // 543
-1.179567765326453e-02, // 544
 1.199294841689739e-02, // 545
 2.696253719652706e-03, // 546
-4.174666056089745e+01, // 547
-8.994533011983796e+00, // 548
 2.471470934375547e+00, // 549
 8.414265353235795e-02, // 550
 1.851569896787947e-04, // 551
 2.825688390924148e+01, // 552
-3.892698665831344e-01, // 553
-3.740765683029019e+01, // 554
-5.173122659775787e-05, // 555
-9.508077249766438e-01, // 556
 2.252008989633557e-01, // 557
-2.657950763992180e-01, // 558
-3.910882557417457e-05, // 559
-1.539077021977990e+00, // 560
 5.096442490053898e-01, // 561
 8.942421981106081e+00, // 562
-3.791455186241816e+01, // 563
-2.210000052710430e+00, // 564
 4.953463876936824e-01, // 565
 1.737931533968977e+01, // 566
 6.530720076069141e-01, // 567
 2.036384610475383e-01, // 568
-1.396017790479317e-02, // 569
 7.116173193188868e+01, // 570
 2.453373197616343e-02, // 571
-8.720524380587192e+01, // 572
 9.547313339820321e-01, // 573
 2.537333920296259e+00, // 574
-7.122460418879970e-02, // 575
 3.749251462325293e-04, // 576
 5.404863282428174e-02, // 577
 4.456197735439298e-01, // 578
-9.676484320706061e+00, // 579
-1.334689593248344e-01, // 580
 1.192766816917028e+01, // 581
 3.750635460509038e+01, // 582
 6.419312208168095e+00, // 583
 3.011655116923769e-01, // 584
-2.329060297931501e-04, // 585
-1.057380976794269e-01, // 586
 1.584016446036522e-03, // 587
-3.815937498960309e+01, // 588
 5.627784116804828e-03, // 589
-1.529300027018790e+01, // 590
 4.313285745235061e+01, // 591
-1.180997907487072e+00, // 592
 9.320946843645449e-01, // 593
-4.762438505497784e+01, // 594
-2.919984874966182e+01, // 595
 4.592501410519752e-02; // 596

}
