netcdf x2b_A1B2Z2_D1E2_v1x {
  // global attributes 
  :name = "x2b_A1B2Z2_D1E2_v1x<3>";
  :d_intra_AB =  2.205224946485184e+00; // A^(-1))
  :k_intra_AB =  7.723480773328080e-02; // A^(-1))
  :d_intra_BB =  1.279961415227759e+00; // A^(-1))
  :k_intra_BB =  5.904419412411548e-02; // A^(-1))
  :d_intra_DE =  2.613944233421457e+00; // A^(-1))
  :k_intra_DE =  7.179196999889030e-01; // A^(-1))
  :d_intra_EE =  2.997713575953103e+00; // A^(-1))
  :k_intra_EE =  7.567530633258577e-01; // A^(-1))
  :d_AD =  1.468342935357421e+00; // A^(-1))
  :k_AD =  8.919884859945887e-01; // A^(-1))
  :d_AE =  3.051790788320679e+00; // A^(-1))
  :k_AE =  1.252270114559383e-01; // A^(-1))
  :d_BD =  1.993046899475141e+00; // A^(-1))
  :k_BD =  2.080854766056480e+00; // A^(-1))
  :d_BE =  2.358253629047993e+00; // A^(-1))
  :k_BE =  2.269127236387784e+00; // A^(-1))
  :d_DZ =  3.702870842776683e+00; // A^(-1))
  :k_DZ =  1.181091190890141e+00; // A^(-1))
  :d_EZ =  3.706169087700505e+00; // A^(-1))
  :k_EZ =  2.861967382715421e+00; // A^(-1))
  :r2i =  6.000000000000000e+00; // A
  :r2f =  7.000000000000000e+00; // A
  dimensions:
  poly = 492;
  variables:
    double poly(poly);
data:
poly =
-3.502242977653890e+02, // 0
 8.237816707425200e+02, // 1
-1.755222230188684e+03, // 2
 2.915862577614449e+02, // 3
 7.557656978745927e+00, // 4
-9.726966146908658e+02, // 5
-5.929698793451181e-04, // 6
 1.176313084884016e+00, // 7
 3.133449537053555e+03, // 8
-6.590624893097595e+02, // 9
 7.388298523020337e+01, // 10
 1.419991332805097e+03, // 11
 7.486617062243093e+02, // 12
-7.315268412498032e+02, // 13
 5.482034399299912e+01, // 14
-7.899635827309351e+02, // 15
-3.608375911898118e+03, // 16
-9.607041798312123e-02, // 17
-1.378998118213888e+00, // 18
-9.187335687306852e+00, // 19
 7.363583968331174e+02, // 20
 9.609524120769167e+02, // 21
 5.765206360617090e+00, // 22
-1.890534095320950e-01, // 23
 1.547884046035385e+01, // 24
-1.455141693418773e+03, // 25
 1.491228756150889e+03, // 26
 5.381848035707810e+00, // 27
-6.595490851879002e-04, // 28
-6.732744432974748e+01, // 29
 9.019616239868176e+01, // 30
 1.086347298021278e+00, // 31
-7.685281461612329e+00, // 32
 5.074825477747091e-03, // 33
 2.431405745835865e+01, // 34
 4.291369336003876e+01, // 35
-4.131352838677343e+02, // 36
 1.765439503185158e+01, // 37
 4.887750470380433e+02, // 38
 1.190131454308617e+02, // 39
-1.044036829655821e+00, // 40
-3.099693347022194e-01, // 41
 4.688086010180954e+00, // 42
 1.072249941975042e+01, // 43
 8.335452670827870e+01, // 44
 1.308140019204779e+02, // 45
 3.565120731521922e+02, // 46
-6.839175005113941e+02, // 47
-1.140863347953583e+03, // 48
 7.431896470902348e+02, // 49
 3.900126803323612e+03, // 50
-2.850768550535507e+00, // 51
-3.319437411357398e+03, // 52
 4.205994410172124e+02, // 53
-5.904130499443309e+02, // 54
 2.111053265049537e-01, // 55
 2.920163463885085e+00, // 56
-3.567984523854615e+02, // 57
-3.492331724067639e+02, // 58
 1.768180115282131e+02, // 59
-3.633657503827122e+02, // 60
-1.457914034729266e+01, // 61
 1.163906366738809e+03, // 62
-5.999720236138188e+00, // 63
-2.177399713514291e-01, // 64
 2.340515068830013e+03, // 65
 4.945830867927126e+02, // 66
-1.863472065745768e+02, // 67
 1.847596401972640e+02, // 68
 7.452808003154017e+01, // 69
 9.561830252494364e-03, // 70
 3.696689935841753e-02, // 71
-2.577869446143539e+00, // 72
-1.946781320496716e-01, // 73
-9.416113634523457e-04, // 74
-7.478941832515537e-02, // 75
-3.858399232268084e-07, // 76
-8.675127475202957e+01, // 77
-5.297675361361416e+01, // 78
-2.955055533113324e-03, // 79
-3.288862550243303e-01, // 80
-8.929466919243973e-05, // 81
-5.863182720996638e-02, // 82
 4.167699151631245e-03, // 83
 2.375885526849007e-03, // 84
-1.907325698645408e-01, // 85
-2.207451676510219e-03, // 86
 5.574876045546721e+02, // 87
 2.723162284564180e+01, // 88
 6.778201932445977e+01, // 89
-5.003723347458452e+00, // 90
-9.040197162061423e+01, // 91
 2.190271928002442e+02, // 92
 4.696131728752836e-01, // 93
 3.949804622582271e+00, // 94
-1.520208939287189e-01, // 95
 3.078608258016834e+01, // 96
-1.319789038049445e+02, // 97
-2.262451298309902e-03, // 98
-1.508378010939087e+02, // 99
-4.950418660917961e+01, // 100
 5.370055859276726e+00, // 101
-7.695504150598895e+02, // 102
 1.722150969638724e+02, // 103
 2.140747104302517e-03, // 104
-1.475962403121194e+02, // 105
 2.672875795070352e+01, // 106
 2.423804438479450e-02, // 107
-1.041699893836516e-03, // 108
 7.616479008302614e-02, // 109
-4.975575096633587e-02, // 110
 1.079033167921072e-02, // 111
 4.603912237507697e-05, // 112
 1.973084765590555e-05, // 113
-8.274918961780904e-03, // 114
 5.562540177071517e-04, // 115
-1.254566578084747e+00, // 116
-3.943003941845976e-02, // 117
-6.561300111481193e-01, // 118
-1.983637136915916e+01, // 119
-1.077760249560745e+03, // 120
-7.324650696518737e-03, // 121
-3.324390272197840e-01, // 122
 2.387671123189170e+01, // 123
-9.113062589386736e-01, // 124
-1.124612450455824e+01, // 125
-6.820402073542676e+00, // 126
 9.876687392375491e+00, // 127
-9.183582067211516e+00, // 128
 1.322628769730215e-01, // 129
 2.257204210881395e+02, // 130
-1.657468591668003e-01, // 131
-7.637940306895709e-01, // 132
 3.941451700845295e+02, // 133
-9.666373940768379e+01, // 134
-4.339415757950836e+02, // 135
 1.408846475323988e-03, // 136
 6.763607796245120e+01, // 137
 7.038607894587321e+01, // 138
 5.208102611197090e-03, // 139
-3.621322384791172e-01, // 140
-1.863788663717596e+01, // 141
 3.136724700714976e+02, // 142
-3.711124899386661e-01, // 143
-1.097551564787192e-04, // 144
 9.445210142831331e-02, // 145
-1.413072525141011e+01, // 146
 2.782289553464190e+01, // 147
 6.642980812291258e-06, // 148
 1.680388122110049e+00, // 149
-4.237634888468604e+01, // 150
 7.955106662990522e+01, // 151
 6.561359551107481e-01, // 152
-4.255819329651114e-05, // 153
-5.895312882458900e-07, // 154
 3.073356469548246e-03, // 155
 2.532315276954287e+00, // 156
 6.415809376259516e+01, // 157
 1.075621245889417e-02, // 158
-4.323576290083677e-03, // 159
-3.611458108829546e+02, // 160
 2.056525309565944e+02, // 161
-9.601964338943075e+00, // 162
 6.682972015312444e+02, // 163
 4.478757398948256e-01, // 164
 1.699133698632456e+00, // 165
-5.687897529570460e+00, // 166
 2.207038488962886e+00, // 167
-4.506007110923275e+02, // 168
-6.491358407679965e+01, // 169
 6.883346963329426e+01, // 170
 2.079260092903086e-01, // 171
-9.349569398563457e+01, // 172
-1.122454304130454e+01, // 173
-2.196727107535716e-05, // 174
-2.573551665509294e-02, // 175
 2.644384779078166e+01, // 176
-9.860420017867693e+00, // 177
 3.272715417085544e-03, // 178
 4.658756664476415e+02, // 179
-7.551872045291424e+00, // 180
-2.743535173714509e+00, // 181
-1.397448928820866e+01, // 182
-4.203227705213351e+01, // 183
-5.963922479552560e+02, // 184
 7.043584211767471e+02, // 185
-1.047485198594917e+01, // 186
 4.136490198818775e-07, // 187
 3.655865044559261e-06, // 188
-2.297390582377239e+02, // 189
 1.981361036693736e-02, // 190
 3.160146247660904e+03, // 191
-1.670138295665171e+00, // 192
 8.717936687499746e+00, // 193
-1.423923426206290e-05, // 194
-5.399508662557636e+00, // 195
 1.244882347859207e-04, // 196
 6.765473887540482e-02, // 197
 2.183776181600594e-04, // 198
-8.407935663504422e-02, // 199
 9.291860200154339e+01, // 200
 1.535591212009040e-05, // 201
-1.396978051553762e+00, // 202
-9.446901131594388e-01, // 203
 4.134642624835058e-04, // 204
 2.219434780794500e+00, // 205
 3.624782985488051e+00, // 206
-6.636828149605910e-01, // 207
 8.782667168388250e-01, // 208
-5.895191713673525e-02, // 209
 6.603585981308800e-02, // 210
-4.819928546570259e+02, // 211
 2.633070802053741e+01, // 212
 2.798190873037443e+00, // 213
-3.016689460319790e-06, // 214
 7.648296782086034e+01, // 215
 1.488148835481150e+01, // 216
-6.399524074993777e+01, // 217
-4.497907080081495e-02, // 218
 1.286976935432359e+01, // 219
 4.038281214321270e+01, // 220
 2.917614069552921e-04, // 221
-6.327687554441943e-07, // 222
-2.021753282298128e+00, // 223
-5.656192607032752e+01, // 224
-1.435491239874497e-01, // 225
-2.051647159380612e-04, // 226
 2.282492479984201e+02, // 227
-1.921839339787553e-03, // 228
-8.146975522560601e+01, // 229
 1.837693869850309e+02, // 230
 1.201084140436720e+02, // 231
 7.364014494468268e-02, // 232
 2.378208562505634e-03, // 233
-1.625310946974404e+01, // 234
 2.259836034811879e+01, // 235
-1.406621282885306e+02, // 236
 1.647420429169120e+02, // 237
 4.613159887074514e+03, // 238
-2.150966625413897e+02, // 239
 1.698876942605793e-03, // 240
 1.159211058436047e-02, // 241
 9.406778870368926e+01, // 242
 1.278939889762248e-04, // 243
 1.764113177471114e-05, // 244
-2.273552240989789e-05, // 245
 3.772964450347972e-02, // 246
 6.351358747006382e-02, // 247
-4.451236136883585e+00, // 248
 7.302710272299662e+00, // 249
 1.041006289760237e+00, // 250
 7.188480849922620e+01, // 251
 5.951954186039067e+00, // 252
 3.914745423828289e+02, // 253
 2.367466745272288e-02, // 254
-4.048521344263569e-02, // 255
 1.113509233050392e-06, // 256
 1.832218659913524e-02, // 257
 9.346654429767751e-01, // 258
 1.072549288071770e+02, // 259
-6.973433452870959e+02, // 260
 4.430029869128251e+01, // 261
-2.118331403818114e+00, // 262
-6.918437887016533e+01, // 263
 2.651025497991994e-03, // 264
 2.086117800035144e+02, // 265
-2.844603552332885e+01, // 266
-2.875662938622638e+00, // 267
 2.891288570673241e+01, // 268
-3.042777771358019e-03, // 269
-2.458942441062095e-07, // 270
 1.015935913909030e+02, // 271
 1.587385041268094e-01, // 272
-1.806160569833384e+01, // 273
 3.262949874076974e-04, // 274
 1.569398068758907e-01, // 275
-6.571050965288806e-03, // 276
 1.956957054799542e-03, // 277
 1.468259388097972e-02, // 278
-1.757779063815011e-01, // 279
-2.649284358402309e-04, // 280
-2.834027565304614e-03, // 281
 3.922180136946607e+02, // 282
 1.030818861036262e+00, // 283
-6.591753621517980e+02, // 284
 9.167604716906321e-05, // 285
 1.345817023738867e+03, // 286
 7.757630650485180e-02, // 287
 1.593291886343163e+00, // 288
 2.404176079938536e-02, // 289
 3.257485300324239e+01, // 290
-6.916828124140337e-01, // 291
-5.710010236653879e+03, // 292
 1.159984584141253e-02, // 293
 1.895463971208865e+03, // 294
 4.010763602466731e+00, // 295
 2.028199176223956e+02, // 296
 1.561381346832187e+00, // 297
 5.541157288810124e-02, // 298
 3.328042453372856e-03, // 299
 1.310449813038242e+01, // 300
 1.298100381260196e-01, // 301
-3.265540429151557e+00, // 302
-3.305796635180602e-04, // 303
 3.517987008693936e+00, // 304
 2.487233779060704e+00, // 305
 3.546762852277422e-03, // 306
-4.571451555820996e+03, // 307
-1.232550365198243e+02, // 308
 3.171573971799355e-01, // 309
 8.046786779440176e-04, // 310
-3.679958458827662e+00, // 311
-7.579349525114678e-03, // 312
 9.785119450527498e+00, // 313
-1.313498475099646e-03, // 314
-4.665830150506566e-02, // 315
-8.494710704861953e+01, // 316
-3.171045384272875e-01, // 317
-1.730016923513933e+01, // 318
 6.258546119193020e-06, // 319
-1.564575182494369e+03, // 320
 1.639731915791309e+02, // 321
 5.104537239747121e-02, // 322
-3.058074166168574e-02, // 323
 1.744781567598951e-01, // 324
 2.589092325893216e-05, // 325
-1.873977175743333e+00, // 326
-1.143105682024369e-01, // 327
 1.522873845329170e+01, // 328
 9.914217017076742e+02, // 329
-5.310536020212583e+02, // 330
-1.284293773927402e-04, // 331
 2.489364470034612e+02, // 332
-1.895181820231673e+01, // 333
 4.442309997792556e-01, // 334
 1.316904858495701e+00, // 335
 2.332480252323809e-02, // 336
 7.332781513117873e-01, // 337
 4.200180758976526e+03, // 338
 5.014934954780814e-04, // 339
 3.929303794898255e+02, // 340
 5.675980977807647e+01, // 341
-1.008441575061774e+02, // 342
-1.123550517718816e+03, // 343
 4.194425719784975e+02, // 344
-8.223879707369375e-01, // 345
-5.890183373523258e+01, // 346
-4.608446584196719e-04, // 347
-8.954922126185313e-03, // 348
-3.294807458565817e+00, // 349
 2.470715302425052e+02, // 350
 1.731911124851557e+03, // 351
-1.235347638508024e-01, // 352
-9.599477266852499e-07, // 353
-2.243501406479996e-04, // 354
 8.030118884486369e-01, // 355
-2.328999127682233e+01, // 356
-7.305196365774883e+00, // 357
 2.167045374295169e-02, // 358
 1.485748204600053e-04, // 359
-6.480085553263185e-01, // 360
 5.175339947173645e-01, // 361
 2.440619553550900e+01, // 362
 5.487563365078989e-03, // 363
 2.346540484885054e+00, // 364
 3.600691876937263e+02, // 365
 6.440814598775918e+00, // 366
 7.380894842768910e+01, // 367
-4.346765990432095e+01, // 368
 1.264933172787824e+02, // 369
 2.059530249240675e+00, // 370
 5.746133019898958e+02, // 371
-4.986889776026056e+01, // 372
 2.889681065479575e+01, // 373
-4.853638726460490e+01, // 374
-4.068560748056834e-10, // 375
 1.328064279778057e+02, // 376
 7.439200773308175e+01, // 377
 1.716341855585365e+02, // 378
 1.313669292190051e+02, // 379
 2.873950655765797e+03, // 380
 3.270898992726629e+02, // 381
-6.686563913189632e+02, // 382
 5.831932783152112e+00, // 383
-1.282499437740182e+02, // 384
-3.131247620068318e+01, // 385
-1.981009311193313e+03, // 386
 6.495273391284599e+01, // 387
-8.838403818168405e-01, // 388
-8.770151418935750e+01, // 389
-3.336696301896005e+03, // 390
 1.809917806926987e+00, // 391
-1.369106778633922e-02, // 392
 2.068183436936862e-02, // 393
 3.143285117391899e-05, // 394
 4.219238962876534e+00, // 395
 2.371702244552663e-02, // 396
 1.005373405361585e+02, // 397
 1.075586896202897e+02, // 398
-1.313150222921167e+02, // 399
-2.492857989702883e-09, // 400
 1.379644394188037e-01, // 401
 5.479216875009734e-01, // 402
 4.587814282796918e+02, // 403
 1.727909208044910e+00, // 404
 4.101384153372356e-01, // 405
-1.770748315541251e-02, // 406
 1.392349684548284e-04, // 407
 1.143829270797483e-01, // 408
-3.488181233167580e+02, // 409
 1.133030696024742e+00, // 410
-3.855495619748863e-01, // 411
 1.507966459877364e+00, // 412
 2.919252998037817e-01, // 413
 4.664698643060618e+01, // 414
-2.725505280626257e-03, // 415
 1.464655388581694e+01, // 416
-4.103921047094330e+01, // 417
-1.748729335502910e-01, // 418
 1.553985899441407e-01, // 419
-1.063701832868571e+01, // 420
-1.276583254474972e+03, // 421
-7.486274994307400e-02, // 422
 7.281615313817762e-02, // 423
-5.269625743466488e-04, // 424
-1.353276657342130e+02, // 425
-8.689124203197784e+02, // 426
-1.889586387744363e-01, // 427
 1.254802125473870e-01, // 428
-8.755040055249630e-01, // 429
-1.150328327815969e+02, // 430
 8.227639828653827e+02, // 431
 4.835092122435975e-01, // 432
-4.206775297082552e+00, // 433
-4.714666649067359e+01, // 434
-8.577684622820321e-02, // 435
-7.601630970931488e+00, // 436
-9.870059105685793e+02, // 437
-5.945767975434038e-05, // 438
-2.293814151631430e+03, // 439
-4.332848397227840e-01, // 440
 1.594884712823623e+02, // 441
 2.101699222796322e+03, // 442
-3.875411721433281e+01, // 443
 1.954945550661418e+00, // 444
-2.751781506644202e-04, // 445
-4.764273534513026e+02, // 446
-1.412486799625107e+03, // 447
 6.489207367084174e-05, // 448
-7.527370359068462e+01, // 449
-8.757897744780357e+01, // 450
-3.634019195049937e-02, // 451
-2.503296726039529e-01, // 452
-1.447162633867024e+00, // 453
 1.891301606272525e+03, // 454
 5.293930903493819e+01, // 455
-3.463540812606311e-04, // 456
 4.576941368363541e+01, // 457
 1.205294788147923e-01, // 458
-1.051840740744586e+02, // 459
-1.888995449415268e+02, // 460
-1.023413822644368e+01, // 461
-5.399332447289993e+02, // 462
-4.335149465073440e+02, // 463
-5.807824600065524e+02, // 464
-4.842381532680595e+02, // 465
-9.437030881683075e+00, // 466
 5.110132681351600e-01, // 467
 4.384760395614641e+01, // 468
-1.023073675286575e+00, // 469
-1.823266889128991e-02, // 470
-8.174997475977017e-02, // 471
-3.071504006898340e+02, // 472
 1.082560807306526e-03, // 473
 2.391201497936088e+02, // 474
 6.232412565293053e+01, // 475
-2.972340660840696e+02, // 476
 4.158550606552312e-06, // 477
 9.829326393823902e+01, // 478
 4.517847153796390e+01, // 479
-7.651894250359970e+00, // 480
-1.143130287774150e+04, // 481
 1.061779209695628e+03, // 482
 1.239626769199500e+02, // 483
-5.293630812167191e+03, // 484
 7.876004728065196e+03, // 485
 2.036781630629758e+00, // 486
 2.924663188599534e+02, // 487
-3.627955559823311e+01, // 488
-3.664823834835784e+03, // 489
 2.661444297514095e-03, // 490
-1.343218817835802e+03; // 491

}
