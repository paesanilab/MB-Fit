netcdf x2b_A1B2Z2_D1E2_v1x {
  // global attributes 
  :name = "x2b_A1B2Z2_D1E2_v1x<3>";
  :d_intra_AB =  4.351828499087061e-01; // A^(-1))
  :k_intra_AB =  7.871036455582375e-01; // A^(-1))
  :d_intra_BB =  6.123463437674427e-01; // A^(-1))
  :k_intra_BB =  1.794150174602620e+00; // A^(-1))
  :d_intra_DE =  2.254999221273738e-01; // A^(-1))
  :k_intra_DE =  5.616209432344719e-01; // A^(-1))
  :d_intra_EE =  2.348979844236523e+00; // A^(-1))
  :k_intra_EE =  1.677719431298343e+00; // A^(-1))
  :d_AD =  2.917299341959079e+00; // A^(-1))
  :k_AD =  2.819793062252046e+00; // A^(-1))
  :d_AE =  2.444010386292637e+00; // A^(-1))
  :k_AE =  2.725353650511642e+00; // A^(-1))
  :d_BD =  4.992136163021810e+00; // A^(-1))
  :k_BD =  2.783935464455248e+00; // A^(-1))
  :d_BE =  2.399566745793650e+00; // A^(-1))
  :k_BE =  1.367713159182524e+00; // A^(-1))
  :d_DZ =  5.972307189645294e-01; // A^(-1))
  :k_DZ =  8.029007089370619e-01; // A^(-1))
  :d_EZ =  1.060879914698631e-01; // A^(-1))
  :k_EZ =  2.311213230050760e+00; // A^(-1))
  :r2i =  6.000000000000000e+00; // A
  :r2f =  7.000000000000000e+00; // A
  dimensions:
  poly = 492;
  variables:
    double poly(poly);
data:
poly =
-1.841049145869009e+00, // 0
 2.596615334624643e+00, // 1
 6.864644234936834e+00, // 2
-1.022900023121498e+00, // 3
-6.702863091072399e+00, // 4
-1.505682788848377e+01, // 5
-3.596680606303750e+00, // 6
-1.101872631332883e+01, // 7
 1.126818700496893e-02, // 8
 4.625956505724206e-02, // 9
-1.083711205651948e-01, // 10
-4.959572652852230e-01, // 11
 2.404993396692557e-01, // 12
 8.650455369211208e+00, // 13
-4.813741745322591e+00, // 14
 2.083395658986073e+00, // 15
-5.183107641760708e-02, // 16
-2.021149768208141e+01, // 17
-1.196040493348427e-01, // 18
-3.098839775992350e-03, // 19
-1.060779419549538e+01, // 20
 2.933482348619863e+00, // 21
-2.471345094666285e-03, // 22
-3.697695277309074e-01, // 23
-2.956368561151158e+00, // 24
-2.103274888541702e+00, // 25
-2.068544173956093e+00, // 26
-2.413557927687789e+00, // 27
 1.874329601922210e+01, // 28
 6.239369718870519e+00, // 29
 6.038034610028249e+00, // 30
 5.283851942097283e-01, // 31
 9.405261094035557e+00, // 32
-1.415665788588929e+00, // 33
 1.353505776920017e+01, // 34
 1.268617293809512e+01, // 35
-3.522680648552872e+00, // 36
-1.022319064418365e-08, // 37
 3.158748035784677e-03, // 38
-5.845963094214677e+00, // 39
-4.271323088558012e+00, // 40
 1.555823829170753e+00, // 41
-7.752831710502197e+00, // 42
-1.183559215099451e+01, // 43
-3.685711088847839e+00, // 44
-5.321108384788426e+00, // 45
-5.860426441813375e+00, // 46
 1.848022862702978e-01, // 47
 1.537689279440162e+00, // 48
-9.503661980547346e+00, // 49
-8.236300035933161e-02, // 50
-2.034681432428248e+00, // 51
 2.370569523900909e-04, // 52
-4.863767101906864e+00, // 53
-2.136342943492953e+00, // 54
 4.543203965062578e+00, // 55
 1.855792193176299e+01, // 56
-6.794687668082750e+00, // 57
-9.883718427816317e+00, // 58
-1.558598698370432e+01, // 59
 3.403068054854200e+00, // 60
 6.495230742293217e+00, // 61
 2.302860363742336e-01, // 62
-6.867507432384747e+00, // 63
-2.334978602326761e+00, // 64
 1.070662663525115e+01, // 65
-3.283244643007305e+00, // 66
 1.480728050140076e+00, // 67
-3.541214401661160e+00, // 68
 6.410215251997505e-07, // 69
-1.971154216549595e+00, // 70
 2.549609140577226e-01, // 71
-5.121524954261982e+00, // 72
-2.298392724346844e+01, // 73
-9.989330692331837e+00, // 74
-2.141385711913117e+01, // 75
 8.493207350713219e-02, // 76
-1.143100399766824e-01, // 77
 1.200075313969343e+01, // 78
-8.837760090724711e-01, // 79
 8.318845529727959e+00, // 80
 2.207448481275218e-02, // 81
 1.414604849208450e+01, // 82
-1.512286862836711e+01, // 83
 1.816781218001065e+00, // 84
 1.462834430750232e+00, // 85
-7.569226188728222e+00, // 86
 9.944998608173672e-05, // 87
 7.256886189708237e-03, // 88
 3.820389017528648e+00, // 89
 9.529056206028265e+00, // 90
-1.913278259779598e+00, // 91
 1.705928831623265e+00, // 92
-8.854235257261143e+00, // 93
-4.287381567454708e-04, // 94
 6.913169460617554e+00, // 95
-3.301318052546126e-01, // 96
-8.758084341092505e-01, // 97
-1.412387932534450e-01, // 98
-1.060057629927713e+00, // 99
-1.935089614520727e+01, // 100
-8.942178544383489e-11, // 101
-2.069962617424366e-06, // 102
-4.483524561888822e-02, // 103
-5.347755592818194e-01, // 104
-1.818037929284687e-02, // 105
-1.286206463428809e+01, // 106
-9.689628253483262e-10, // 107
 1.605783294772072e+01, // 108
-1.230878743953684e-03, // 109
-6.087492932149734e-04, // 110
-7.189246640339252e-02, // 111
 7.512083896475442e+00, // 112
-3.958296085974248e+00, // 113
-1.438752940957272e+00, // 114
 6.312543804244256e+00, // 115
-9.483859815781809e-02, // 116
-1.466417106112931e+01, // 117
-8.467820489824886e+00, // 118
-8.733738865702980e-04, // 119
-3.826197696821190e-04, // 120
 4.976124665226301e-05, // 121
-2.160799547240840e-04, // 122
 1.413040829830447e-03, // 123
-6.128738262423088e-02, // 124
-6.959820684523961e-05, // 125
-9.702060662574045e+00, // 126
-1.500105072178108e+00, // 127
-3.309466819081639e-08, // 128
 2.611133712025009e+00, // 129
-1.630866772082432e-01, // 130
 1.125938815309400e+01, // 131
-8.238708959472293e+00, // 132
 2.028140495624237e-01, // 133
-2.751411571564938e+00, // 134
 1.129424768088241e+00, // 135
-2.871940113821929e+00, // 136
 8.052598957423832e+00, // 137
 1.375877965482709e+01, // 138
-3.293933405800950e+00, // 139
-3.733944195060344e+00, // 140
-1.568064213815975e-05, // 141
-2.665979379570448e-05, // 142
 1.473756225675794e-02, // 143
 2.704598790534578e-08, // 144
 1.188666745407006e+00, // 145
 4.062685351651391e-01, // 146
 9.799232144624272e+00, // 147
-1.441477068808277e+01, // 148
 1.802261421595024e-03, // 149
-3.143088825595380e+00, // 150
 1.327616772404295e+01, // 151
-5.510406838647582e-02, // 152
-1.112207607376136e+01, // 153
-1.345924296813404e+01, // 154
-1.424691642803437e+01, // 155
 9.421550842980199e+00, // 156
 7.217455327926174e+00, // 157
 4.254244969521210e+00, // 158
-8.611915387176118e+00, // 159
-3.408866200493472e-03, // 160
 4.208097081074345e+00, // 161
-9.269178930942350e-05, // 162
-1.239011324526440e-03, // 163
-1.867711189786185e+01, // 164
 8.833546667591869e-04, // 165
-1.000684428154562e-01, // 166
-2.220881244223389e+00, // 167
 5.073865875992876e-01, // 168
-1.394516754837034e+01, // 169
 3.349550549060920e+00, // 170
 3.338038350053310e+00, // 171
-9.338294615088841e-03, // 172
 4.685674338295483e+00, // 173
-7.852422619763772e+00, // 174
 4.261436558150246e-02, // 175
-5.286995544063805e-01, // 176
-1.836992470754056e-09, // 177
 4.847490206758891e-05, // 178
 3.335498216756393e-06, // 179
-6.137069309638063e-02, // 180
-6.307780873582735e+00, // 181
 6.948630622298499e-02, // 182
-2.917335977911817e+00, // 183
 2.081316616422872e-03, // 184
 6.915316427580338e-04, // 185
 2.830786341810249e-01, // 186
 7.968011347705414e+00, // 187
 3.002972954199114e+01, // 188
-1.072547209998409e-05, // 189
 9.641806694417788e-01, // 190
-1.197398805170560e-04, // 191
 1.345252492058653e+01, // 192
 9.860900031711331e+00, // 193
-5.965304652693291e+00, // 194
-1.883132003642447e+01, // 195
 2.527024285182730e-03, // 196
-9.286948738376756e-01, // 197
-1.897399016085030e-03, // 198
 7.340930698424908e+00, // 199
 8.579308106116974e+00, // 200
-2.262448363749524e+00, // 201
 7.566230174112491e-04, // 202
 9.119399927301369e-02, // 203
-5.698140975922788e+00, // 204
-1.150712536825071e+01, // 205
 6.689066193822519e+00, // 206
 8.931125209671200e-01, // 207
-4.382606910945016e+00, // 208
 2.116885686626013e+00, // 209
-1.009318463885531e-08, // 210
 6.492602473352045e-02, // 211
-1.224503564439979e+01, // 212
-4.755212090461615e-01, // 213
 6.398431031065863e-02, // 214
 7.919863309411841e-03, // 215
 1.523205152026107e-06, // 216
-2.189880951565548e-07, // 217
 9.210381529462706e-02, // 218
-1.069762662481852e+00, // 219
 5.563358660146127e+00, // 220
-9.408242547284443e+00, // 221
-3.224435391612661e+00, // 222
-2.399766313351115e-04, // 223
-3.184482505634387e-01, // 224
-4.948153891962180e+00, // 225
-1.376312076211219e+00, // 226
-5.204474967738005e+00, // 227
 1.958990924982251e+00, // 228
-9.877904136069329e-01, // 229
-2.690388224308824e+00, // 230
 3.266631556969330e-01, // 231
-4.825587489196360e-01, // 232
-4.724630758986102e+00, // 233
-3.340078307978356e+00, // 234
-1.783909928084840e+00, // 235
-6.689974557106653e+00, // 236
 2.402263644525786e-01, // 237
-4.820246067408818e+00, // 238
 1.441771077966689e+01, // 239
-1.019148948131067e+00, // 240
 1.541171360790910e+01, // 241
-7.394352323521792e+00, // 242
 5.852572004179975e+00, // 243
 9.161709371005734e-04, // 244
-2.142835592809065e+01, // 245
 7.073849212318460e+00, // 246
-5.835449823534172e+00, // 247
 2.013144585531750e-01, // 248
 1.305940471326016e+01, // 249
 2.618493280993485e-04, // 250
-7.908405327290970e-04, // 251
-3.753752380084114e+00, // 252
-1.165194396885548e+01, // 253
 6.482231857929071e+00, // 254
-6.781952815076072e+00, // 255
 3.477554879427032e+00, // 256
 6.275920021983841e-02, // 257
-9.976154421045882e+00, // 258
-9.574933726845861e+00, // 259
 1.204270044148915e+01, // 260
-4.273134183470188e+00, // 261
-4.157271829659242e+00, // 262
 2.396133812163992e+00, // 263
 6.547062703611227e-02, // 264
-1.087550418078889e+01, // 265
 9.965988437218909e+00, // 266
 8.142965004081057e-02, // 267
-1.320089554384385e-09, // 268
 2.653091236520382e-01, // 269
-9.363440398209567e-01, // 270
 3.304767110901934e-01, // 271
-2.528596166421435e+00, // 272
 1.117373623195679e+01, // 273
 5.426045159415987e+00, // 274
-7.470695903362989e-04, // 275
 4.040622123210828e-01, // 276
 7.091974935764717e-01, // 277
-2.688313356393402e+01, // 278
-1.752839589952883e+00, // 279
-3.631085256539185e-02, // 280
-2.828459835703503e+00, // 281
 6.780816495498937e-01, // 282
 1.777809893317599e+01, // 283
 1.309174653088738e+00, // 284
 2.490579232931438e+00, // 285
-1.226161510534070e+00, // 286
 1.329407563496377e+01, // 287
 1.438245999113643e-01, // 288
-2.680697326039672e-02, // 289
-9.633842467592014e+00, // 290
 3.092960471703948e+00, // 291
-1.335104191397555e-01, // 292
 6.172035587506343e+00, // 293
-1.638633063213263e-01, // 294
-7.445379289914439e+00, // 295
 6.059958603871145e-02, // 296
 2.341757791840375e+01, // 297
-1.052761117215334e+01, // 298
-8.304478774969315e+00, // 299
 5.910179042230760e-04, // 300
-6.580040858324666e+00, // 301
-4.625911243618230e+00, // 302
 8.460719375580604e+00, // 303
 1.185347701565721e-02, // 304
 2.153194635979308e+00, // 305
 2.496177509686474e-01, // 306
-4.737468619814880e-02, // 307
 1.914575862118107e+01, // 308
 7.434271227529126e-01, // 309
 1.711479091489334e+01, // 310
 2.847268585064802e+01, // 311
 6.925265808390804e+00, // 312
-4.643061379138285e+00, // 313
-1.964991819100593e+00, // 314
 2.861403610408022e+00, // 315
 4.822306119584529e+00, // 316
 9.931182457918280e-03, // 317
 2.462223620367669e+01, // 318
-5.242463962011088e+00, // 319
 1.269988752473649e-01, // 320
-2.791246058864554e-01, // 321
 3.439090329656157e+00, // 322
-9.921042466663147e-01, // 323
-1.193400958282707e+01, // 324
 1.691560429504198e+01, // 325
 2.659432551680709e-08, // 326
-1.028471700106001e-05, // 327
 3.890261170127605e-04, // 328
 1.483715573392777e-02, // 329
 1.075710473540759e+01, // 330
 4.802678355406483e+00, // 331
 2.137766688230261e-07, // 332
-2.072535809601634e-02, // 333
-1.699050322952613e+01, // 334
 3.909281439247505e+00, // 335
 5.862416077764513e+00, // 336
-2.301976850682115e-07, // 337
 1.348568156138561e-03, // 338
-8.298679853432066e+00, // 339
 1.551481910735483e+01, // 340
-2.706085295927768e+00, // 341
-3.145855502190065e+00, // 342
-8.981319271076597e-05, // 343
 1.092166058577906e+01, // 344
 1.291746470046646e+01, // 345
-3.497495927975645e-01, // 346
 1.085823920119067e+01, // 347
 1.602623994667150e-04, // 348
-9.512539813169767e-04, // 349
-6.184161252832530e+00, // 350
 2.484983861033316e-02, // 351
-1.514824556983484e+00, // 352
 6.095183230085664e+00, // 353
 1.033412781514268e+00, // 354
 1.187672369802302e+00, // 355
-4.521540661772163e+00, // 356
-6.820062973110262e-02, // 357
-2.693770707592605e+00, // 358
-1.238987734424573e-06, // 359
-3.994580427077225e+00, // 360
 6.351751818726561e+00, // 361
 7.598306345472558e-09, // 362
-9.162873315653490e-02, // 363
-1.359945106314553e-08, // 364
 9.337742511762462e+00, // 365
-1.337536645973756e+01, // 366
 4.624203232169138e-04, // 367
 4.534410268042732e-03, // 368
-6.801585292256685e-03, // 369
 5.188964429445642e+00, // 370
-7.113272958875989e-05, // 371
-3.032347168427777e+00, // 372
 1.584817855465320e-07, // 373
-6.546913693795555e-01, // 374
-1.082965391230716e+01, // 375
 6.828643309749519e+00, // 376
 4.914748877821945e+00, // 377
-1.395939795212554e+01, // 378
 1.566236166264581e+00, // 379
-1.713912732016619e+01, // 380
-2.068557732135928e+00, // 381
-9.825551785312810e-03, // 382
-3.239243081216433e-03, // 383
-4.025334319523119e+00, // 384
-6.234092655292949e+00, // 385
 2.374004117720913e+01, // 386
 9.757745450152633e+00, // 387
 3.503489501825313e-07, // 388
-9.107510787510606e+00, // 389
 1.631819876427032e-02, // 390
-8.881700685689058e-01, // 391
-1.042117391705776e-10, // 392
-5.958918642861936e-01, // 393
 2.875287598390909e+00, // 394
-7.888870711887372e-02, // 395
 8.547402481975884e-14, // 396
 1.366545961608151e+01, // 397
 5.220467115668957e+00, // 398
-5.650940854732273e+00, // 399
-9.074015207299956e+00, // 400
-1.478393938914094e+00, // 401
 8.223392671783577e+00, // 402
 7.234004243200333e+00, // 403
-1.134543108185613e+01, // 404
-8.307418982717987e+00, // 405
 2.999790860821575e+00, // 406
 3.649193595678747e+00, // 407
 1.216881269445658e+01, // 408
-2.414806773345227e-03, // 409
 1.828582363529319e-06, // 410
 8.751578958969611e-02, // 411
-1.043659686041376e+01, // 412
-1.857064030644103e+01, // 413
-5.228158484627803e-02, // 414
-1.242347518288548e+01, // 415
 1.197707971172004e-07, // 416
 1.032915668662468e-01, // 417
-3.537546268445870e+00, // 418
 1.364716826482437e-03, // 419
-4.848197392311206e-07, // 420
-3.443738631347529e-03, // 421
 2.280497427608200e-04, // 422
 4.755562814871550e+00, // 423
 6.314738767967592e-05, // 424
 4.556442423380497e+00, // 425
 5.319166258360929e+00, // 426
 3.474415406549122e-05, // 427
 3.687836526004355e-08, // 428
 3.239729973944360e-09, // 429
 5.295750554637005e+00, // 430
 2.517819254997451e-02, // 431
 1.202531628109741e+01, // 432
-8.743933024131514e-02, // 433
-5.748859732648691e+00, // 434
-3.216403326937080e+00, // 435
 1.138545219016921e+00, // 436
-8.383271409772554e+00, // 437
 1.615616507850513e+01, // 438
 2.161979782440900e+00, // 439
 1.149631590097323e+01, // 440
-1.041153203140474e+00, // 441
-4.436430841582324e-01, // 442
-2.441264502304078e+00, // 443
 2.396743411430435e-03, // 444
 4.336369381857595e+00, // 445
-1.805523775329794e+00, // 446
 8.111733169485939e-03, // 447
-3.910674656789363e+00, // 448
 2.672629152245604e-02, // 449
-2.464639929994058e+00, // 450
-5.740623107436193e+00, // 451
-4.791286516067002e+00, // 452
 3.611560444112498e+01, // 453
-8.592540261211582e-04, // 454
 1.164679023711054e+01, // 455
 2.969633510655160e+00, // 456
-3.992990313660869e-02, // 457
 2.761710753374968e-14, // 458
-3.672895606601431e+00, // 459
 8.793781050401236e-02, // 460
 2.288362846791640e+00, // 461
-4.536085043809699e-01, // 462
-9.972098212889668e-03, // 463
-4.811939506256093e+00, // 464
 3.218118675005603e-02, // 465
-6.071266851176391e+00, // 466
 3.739226049165599e-02, // 467
 3.104187909419678e-04, // 468
-1.146765716589588e-01, // 469
 6.930951991947870e-05, // 470
-6.682587418849949e+00, // 471
 6.022502943781850e-02, // 472
 1.092519548349924e+01, // 473
 3.500136761841146e-01, // 474
-1.486066171325782e-02, // 475
-3.347429835196309e-03, // 476
-2.152797143100686e-03, // 477
 1.019098048841654e+00, // 478
-3.365738542310761e+00, // 479
-1.615193204093934e-10, // 480
 1.475820548182271e-05, // 481
-2.366384461061946e+00, // 482
 1.249451862630125e+00, // 483
-1.786734148614248e-03, // 484
 1.731838905832005e-03, // 485
 3.863314212966233e+00, // 486
-6.493304876111941e-02, // 487
-3.333794717573472e+00, // 488
 3.415457063896087e+00, // 489
 9.557563116659100e+00, // 490
 8.200324961280064e-02; // 491

}
